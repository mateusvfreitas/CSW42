`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
zEaqTwG8RX4WDqFsN2A8rZGru307yGQ9cgJJdQp6wcIn4Y9PGY8joj+I6xsGQxqM
ZLxrAQKhkoExRrIk5w3qaWYzuuZns9vlnLw1xqDrVcd9lO6FOVM2/UPxu1Xi005D
qyjNOE3hYZlWlrzLZ8MCVCN5p1XKqvwJHWtcU3j1QDb4t+AyioJZUtGtAB3bj5uM
twH3n+tGytDLGIAhdD0we06Izif29n4CC70Dw010nikydJUrj2+8HzIvZlP5XhMq
XC/r8PNRylynNt+27HD5NVLq00KuEW9iGqTrODT+9PnLo9NGQd8DwtTuUVSC4zgF
2Lw2y1kcR9d5PGzH3+B+TFKP+ypsFX89QsDewAzadu0i6rMf3dgjxNwXsl4Q87lK
72g0FW2xRmAX9bNBN3P0WBLn4xk6vMQbYovGpulHWq+xkhWf1hOZxy9oHxajDuWa
0/iIceqBj6Gt0UHmDwmA8YP1hmgrLEDtweUj8hR2UGBgldGwlJUdV76sX03eyGNe
iVIrcoi+4db3qTKHo4G51cChe6sfXU1xFMZQsOd+IAW61VHgR1WBxV8C9aMkZLdX
YUstStZxEqMm/l6+4kmtzvbbbK9Nay6E0e6qVzSwWwcXgLALJ6Y0nJprd5QqMit+
VJ2FUcCU8S6Cje0VdS66M+u1PQZM2aw1H6c+livoFZ147ZmWg0TEq+V8p4250MQ3
zKEsP9P5hhdQKeSFGk7k6GNCC32J72Yk+NDlls5W5YE=
`protect END_PROTECTED
