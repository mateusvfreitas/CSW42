`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ta9oafV5Nlc9WyX1fuoaYk/vdeW0w8tUuop4YKhIYIUqY0eg91IUJQnfyedZ8zT8
Jol0FZ3L6S5+a++2mw59H+eqvX/XmILCByrnrJf27AEsYcqChGMhTLdERMC11naw
80v9saTF4OIagYC9ub4LGWYijfwMVwODM1IMl6Jl4Bvqur8/eQ0rfL90pr5aa+Qt
QozJCzV9GtZSx2fDJSop0WBLh0utP7N4OYeEB1h0HunExZ88juNsZi/ahuhKONYL
sthVujdT5ICzukdmfLYNLvT49K6fqFYfvP8Vl/eTfhPqvOI4zPgRjUcH4uEe1ekV
OHQzEDxzrFlamwwZQqiBvOFp4QKbp6lUEdEm1UbAo3EdHm5p3ZLCrywCeky5nWpF
yjvgNn5GDrsBIyPp0fwc6ZfSG/9dcGEjQF35BM0X81lXVWCXhZfh4lwsP8jptQ0+
Jw5ooYhLjzPQ0G0uaq2RqQQCEDYwzYGkyEOb1SL1uH8KCjaIIAPqJVKFrqQ3Z+5b
HSPeA2vY4a5hAiveMMYCS6mElx8amJHaxHUoaBQkNiSV2Y/tFFaGYsl7hMKcf5Fd
C1Xy84BBqMOeFaoetrDDnSg2U/ojwPhp1eiWYJ1guARvlxr2kqijUco4bqSTTyIm
X/IcD5CS8SH8wtx5/8ni6536P81jfH0IjGfJr7wTBu7wRhLz7CWGHNkdiv3QUm9Y
qLK6dtJyfO0jkhupm0w6XS4Dt4+YPyViEczCY5t3eVgQyYW2qJnymUHEZcuxE93P
R820HqOnKJGgdlnpoNmcbmt8OUDWO2w6dAa1iqUzsdwEz6ehni2C6gEmlvBCo+X7
/4YWC3/3DE9HUiq0qrg1AOALMO7TA1bfJj5p78kBf8I5zgOl8nnDO370ywamlZP4
wqt7puyznSNgK3avN+sxTbSrV5WIwTLLxrtvNKnqge1WFvkBOVMsB55MHH9rfj4D
ItaFd9OkYNPFoAiuQ+XhCoEI4IVXsYK/HBSEcIydocGktcPYGxwUY3pd8J7GaAOd
oraRtC/GzxDYyLtietsV56IeoMJZ8/quil0uiKROCs7NVXxj3dlbEgrJSjthfNOz
uwH2Si19S1+zRSuPY06uJK7IIufBdVrq9xI/OqOP0XdPVT/nn8odyjQV9TuktAxo
ftarV/DR5EQs3DUkrY8rEsjWzwFxxZTw8iM7pDOLBgRfVix4Cd5G+zfI56kbX97m
xCj3fTyXjKykuOazIm4YmsagHt5+V2c1AEDbYAC2lsYByci4KGJizhDZsOtXQGSB
Ojvx7642KMmihu/XHaunmH/PFk/KRUusYpdYtKavBo2u5nfFoGWvuFct0ocUnNTq
Ea1Lil/Hjbb4/w/U7qhUIAS//DAH4Pq5x44FFr4HvN9Vao5BVIOFxdVJxSPdM5wc
BsCTYaZ6oniyQEVOgC7yhrikUViMNC1q5951WEZCyufS1E+wdtaqi4XPII8SuPkF
41JTuWL4E3onh3TUbRWwVmhLaNg0xqhLIr7VxFs/r6AMNgNxvprciu5lq/Bt8/H9
IndS0LYiSSkAYffhxaLuZBa9H+NriqyfseK4jFjSDn2fSJGoK+CcD9TSlkOCN/TC
hapY2PHLWZlndix2V6NADyf9XnYeGvQTS5C3OsW4TNBZQeh0H3nS+8jIxIBTEvWD
D0iQ7X1Wc4rAezC470wmqiexDrtMm1F2jbqqQyZdwVVQ39bKVmHls56rrVRPA5i/
gyQ25vWzF+M2efRI8fUgbMozK0Dt4kqeGCGBuOcQkTihwkEs+TwP87iJQC4nuB5w
6K/F7Q/UwVctfPugpwPasT7keHBqQxNL6m8dIBFeWrk0iond8DpiOppNtqg5yLKo
SWX2sMVKqeri+G5QRwKzVlVekZG8jFvIqH24iaiVGDds6aHYSNBlA8ixdEp9z7ln
Hwh+oxdZTyRkggfTpdALtgHa5Kfzikbz6lhC261jFOOtz8XGKFaSBxvPaeTtcF6R
y77cJbumfWbSvhBs03hlX3etPeC1OwXBGFPv0iyajzDFQZPPh/xjRXfMgx10i+Mc
LZF3aI3B2iLMx6famfTF+w2IneJTZ4QiChqdlyNi+Nri/rd7xA/PMqgog1Zop+QG
BQG9kPMYLvYVCfLC7TqDebViJKOeZrCxhUasf58bXkMkE1vvxmSrHBAk2QxpAO/q
NsDF5V1v1qAWhxKSsznUiRbn5CNpFo5ALrtKPsQp8Wdkow2lEw51GTN4JzQtJhss
0oSvfW/s/pv6NyDVDWSo2Oe0XOAVJ/8MZO/eK3mcTkrrXGDO618L/C1ckVtw4UH1
te+Nh8g0OtJEInVfhWjX4+y+RtposSXGpl+81xk9zF1X1hY2bgo/2b6w/bGAJI8b
cWiSWdRxQ4aPKrgPnZnZVfi9tV1EsA3TsgDQySC1256/LFaloEWB56L8B1U4Vp7s
61S88dCDvN0aexOYrqlYkekdIkGglqwOkoHdMf1AAzarUMsPQw3oWtCFfmqJA/li
SKJeJ9y72sTGRSv3zXxw8qQfdEXmWTCtmgXFGWFwzao32w4v1kCJNarwylZNahi3
GtlI8GQCEChfr4yz3UZIDWkRSW3VdV3R1+QCPTT4uyBfIHqNpHM8nEFBFGkA+15Z
Ekr0QS0XFZAt4vNulKXc5xJQuNCQeR07QfwRMd73nl0bjK0CuzM5yYkwDFqlDkMG
Qgde2qCANf0g84dXySPpsuGgvL+o801JQ/36FAIdtUZ6sfLgdld7tywjs4Hn8mI2
IIk/aS3iiTc1zN3LjprhaFr4PhRdm2n1TCivSQ4LfEKxLkXVXmOFQtbQ2B17xRrF
PTrpStVMQCNoUP0Pjd7Q41sId8vOVLTUZ2+WEYdl4Wpnm76z0Hw4a1cRfrDUYqpc
LothTRE+0/WfW/PZr/BmIEpzH4fHY8n4i494S9da3xEV8GWZYwUY99kAsi+OAfNp
LkezqN79WeNuhjhWE6CCnxZcWAjao4vjzLOQViJKSzNUnpAzlFhh+/Pe2Zxu+GdQ
EhTbQo5VTCMwzqK+Qo7GGCFWBEBEFXGicAmPgTG1SxhwFch3q1GwXGYbpXyXEvr2
EFyFxG+9q+KzROTCrgVtvviMboyMqH89OtnCWkK6l1peCEw1XAVOxw5zCX5lTvsC
qYOG69wKeSY1WfQmM5oPixIgmn/abiUEckhc6asBQmuLCRs2MMdcus3wYtai5KBm
6ZXrSfIdYp27QrhltGqIBhnRBLEEoAHFBf67T3AKEQB3/zZdfL4BhAnX+ygnI+ol
CzSQ5QL/FQNbYUljmZhMAdClA+yeBhsWsOlkaIPCXw35dOORXTwcPMXc4VqNg3Tk
x4J1OfPXniwUSBNqnWS7AyNtcz3G8fzVu4yORPDrxU2dXSAbKANcYiwg16pXPVux
cK2fSo0Onbkgwe3EWJig0b/QBqlKzkdhJ5xrYMY/f7cfvDS6hoDX1MDJmXJpItZc
0Y3NrmanFaRvf5J5uyM4SCOX7ENugvh0DAh7JOf1jerAas6goAwbiNLwUF2n21zi
piGD21iji27p904KErktI1FJFR+y2E68If/mPncQ3ZW831wtZdN1DcTC3wvYaGdj
3Ibw6sdc1RlzBqVD9Y62Ff2AEjRLwAibj83rlMdDIYbYZSKj8foI4EnGHZkKY4U+
iP8Z8Op89qhn7te//TQ5Gdue6oIx1qp3bvCAx17bDzAmYdDrYulb5Lx52t0IwIsw
hRNLxosLtUpaa1s/dzDl7DhxgnTl3rDeBVG0vSqto9yTL4FHuZlUDa3Y6h6KPS8r
hykiI43njpDffyE9KINZ8G3suiaImt9kq/enxk10CQ0MjdJ1IoiyopV8A3u2dBvc
fZ9eCp+nYdUqpeCsn0JW5OzFulssZMrymTWuTK4lXh0pqHwP7layZj9CRqm/PYsy
9dzD1x5ZpqBxRR6Y19gr38nfgAaMhfwrzRc3F8ZKv3w1tcQrNVvS+SGwrLyxBEl2
ZKd/Sw9+OPhkaIc+6upLJkY3XidsBkTwbIlaAqKmistaavKgR8iLD3EAby4zceGN
0YYDdxOdOSoCv8OtUxdn7PaEE+pnbYtHlsQso/NPrEDKy81oVJV/uX1KIM/qCFI/
IgKnDa01DaOHgfh5PUbGltZ6gk4ZiTKWBxiFHAavg3RVSsAz4MiMT/vNYutysKu1
NSTqTdoxenEJYpZpvSjP60A5n1smOd1kUR35P/Rb6GKWHIxvgOGMgISBHnl24wJs
+jtLPOLuKFpkb1H6u2Isw2F1ESwS+eN/SegQ2ZxeXB/P5UGFmfFdqjIUWBQBljMA
ousFofFTY9CAP4YnhrnoLKmqPb3UwvTM7e4OxecFwxCLjDEtgZRNBG9dt0UnIvql
LpCpKlUS3OfOIkWHEbJy1I/13e/MfJuuVU0Uh/oI757onzp3b/EHjnXgwKtFsR+i
lFdGUOCGAuVo6pbKUd5hh9drz9DMRRTdDcOsnUY0bX5oHzjJssAkM3ta5cRmq4o+
p9IEQlyHlS+sQnmbjIJl6hEGJFaR9DjFW1x/7l3QDOlerPXLrfn62fU8W+4Rhc0c
/uO84Tyb023mpThoCFhvh8PyUsmhLQ+yYgRK5kWv3VIytpwOSEUeKPcA7RDyYU9T
7Q/K0RIPBo+QLgPnpze6SDxm/lR5vWK+sNHJHs10bwIUA5fW2mAbO6qoPes3kQbC
4AJfMnz/0fR/L5A0AFZl68K5IBGg2gn7l0tka5N5FQItIEnCLVRkE3juHw40i0rl
V0ZniVFTk6yWDna74i9+Ua+50V8fikuRXDepTXZUQ7a2HV2xLKGc6DN8aqvLiVJM
2XpIpw4L2j8QcW+EKLIbriLQXbODoeSYoiMp+g0Z1nYiq2KBW6Zi6ZeivAIv81J1
UCgLVlDu5F2oHgh8LxGoOQW0Mtl8n/nUwDP9FP8H8ioJyX/Csi91ebBUZrL+bpUC
8FRxaYnKGC/WpkZkcBJ1JAA8EW8/M0oRZqkpKTsWS54/g7llHUm2sBQV9onMEHDl
hzjzfKcYQMazw7XLUkGS9Uwd0v3p42D2LrLsildyzET6ztnLv64NOWtNUvrt5yI+
2oXWuRkoTwCFs5DEkrW/HjixVCuMu+S+wExc+lZnynNGzAKgEIQ9/oS7VZwwGERO
QeLU6Rk4bsKxdyrf3eIS4J05H63Z7xLBTRp4CpXGc+oggl3iSXiqWnWL9FXIu8VL
9VDf9wF+k4P+Pg1zM6ZYgOmaYBQ/IfeX3GAJCC5KiC5SBdMragN9bBM5Sjn89A/J
8TlbVD6hmnh4f70moGBdbJoq6Fb9uhZzUIG/miyVZhZ1Rbrl0zQ87Azry+T9GwdA
insUwwAK9LnnZV5/cwqCzEDQ/Jl5yq1R+es33RuCe7ExbubDBRibfb8eFjw7ZvWM
f5277oA2xHUGHAElVjlOMgst6wLeWRqDbj9KO0t/I7b74Kc95fpv/00dEiNpUNhF
c1whynUagRzPncqHVD4rjndpCu2ekiEJhzBRzAmXilfocuKIrB7p8qt7U/U2bK+k
e+WwRP9lvyJhz6D/HiK0dOHl1hj/63rEkDOFwJrs6JEr8d/TAzyuu14QB7hkPKrG
SQ0IT7+QtffxaE18TkxSfxF2lmx4yyTtSTR0zBVHNYEH/VbbIrgGdvlpudGrDnQZ
IeNCnaPCR3QJWwefg8Ld9RuK5fkzxvXzxihUvzynIw7EBRftBcBa12yKMrzZYMfB
iAC3v0BDDIDW+96idbJObhOC5TK4D/xQxXWxaejVltwCQoer+JezGQ3vsim3dhLQ
dRc3lHywmtBInnGV5jYAqxCFVtVjJXJ+ZMdyRsRM6JuWAV2Di1jQruSbqSVFjdBK
BiDDFwS9qZ9C25qOxSeLCkx73EbozVXqtaHc2lqrxCjQc0TQJNBImjgifhaZw8QF
9+R+ZBORSZ8qP3KP6H8Miip6jStD3kgopQwAaZxedH6dyMhS5+oXno0OrqWwJ1Gk
q/EegDjbpdaWtUnrTLRO+WehaETAELqnsgnjD55+IfMU7T6KOLXh76NU/YbrCV9Y
hFLC7+ApjOpdtZqnLB4cI6mjnm2OY63TMLiUKSYnHiO8flIUBwxUiYiyyyVLMVYn
LLpxdjX6Wp+HtmEjX7a8udXRQP8ID2kNAtj5ZwQtCEUpD4AEurwrjcXjf2RiaocG
gPseXrddouV1nAaFixCjqHK7Ii8b2F09LPmzGawXYFcurYJ5kO71iLE87E3sEAgX
847GRJ6uY3/T0P3WrtCmBJWeUMShy4A7W9EAuMeAt1CZ1x943nP0Ax2aFt6AdIiz
q2oTaihYfaqWOmghL3M+WKf2I2DqdehquVmmYFjK7Txf2frWTOvmMVadrtvXSErv
wOX2bGDc9PmoFMFGLO6U9NxzEwUOY7kvVJdNGPELlnOH87ml4UHN0XWzdFnOJwTE
wfQaUG+z9kF+NTR874ZrUY6ENBL8PTpTkXencdV32wRAzQQ0ML9d97Xx3IhkiSBd
+ViFtMVWhOQmtY2XxjJeEGwLbV/3Nuzh+ZojJQgmvTSA1YmgbOk/5orhv/vvvNrF
AoLyxgleClb4qf4luhBHPY/KMnkln2WDOYiJKL4uPk1PuG4oOF7biXQEZercV3kW
4z27sO9ph/7PlWG7Yys/anDXynklBw7X0L2gotwz77M+NXLNp9STnkMo5yOn+srl
GxRBnFguPvitR2o7fJafc2S27nD6EPd7pdFCVLrwNFjKiatmZdXMBMiOeis3ava9
303SieZ7QaPUFPsVrRHu+L2dLMEL6LRWLZnfJ9d5x6JrQPPxl9mJg7iFm+HKY/ky
LdaojqriTo6fFXElhTxL0nMlcfWpxKUf7nvNrR6t+YKI9XDLruE0xp291JjshTJt
Af+8TvTLXXj4fujCWheWknYhZYU9J13o08zV4X/EAR/Hzm6JpSzSKcPyh6HiviR/
3yS/kO78X18j/ouWJv1HL6xbkqCn9Ua+qLs5TRQZHjZtYWCL4pGjnSYlBR3RRTFO
rg4ZUgvY1SIH0sC5JdCFWRis1RYt+5lD3RDkARkbryTPgMm2VnzEAteLl/f5e9sK
AGBEZNjdLLP/DtnmyUiE5TI5ox26DLxlKfT4qJ5fNChe6/SABq6nZHP/nQ+WWc5a
hhBowii2jiojBFC8dW8OyX4ipgeMWUs/nSKQn/j7xqD7nUtYkE8sDIy19itPW/IA
zWaMLkH7aImr0bIbrfyN4qqcCenK0YxpVettJQQfpZsBiM1FQHAmAfo2NCoKeihO
MZR9iARKYgl0wqnHKghT8klXsOvlsXpmic3UtYtCyJEZf5t+GUMpN+VuiZzqmuef
3OYMMrD0ms+BPORBgOVg6WWHPjIHGsZQqiZrm+p/YQ1BNfBnpi2CazP7nsBXa6gR
t9gMTQegcnb5l6wxZ6ntxLAO4me4zU21cEB1OsxZ3mTXS4tDo3vP1v35lW/iow1B
GdomZ59byy4BH0NhfkPAYJoacM6k6/yUp9KVOPFqIBTK+KdMosnBoMqTalP68Ilm
K4lbgyBme3Os1bjCsaHo/sG6/TOOkLVu5Nc+5YZDAaB2Hgjd5n7hcwxlvX8EniNB
DhRmvpBX3HY4kJZYHtE7u4O+KPDLU+gIhWm/YgNkfgQXAdCrFwqmydLpEXfzkZuE
JD1abEqhYHgetcRfwfeuv8Mnfg7ZDPTCwwqS5D6u/QTuUtJH3yPy3+hiz17qtFlK
6oeJPm5bXNrrHAjSqL8FNSjzU2m028j68+IbXY/RP/L6DwxKN96nTmzuA0QrYdwQ
AcMEgjUeF94sxomFKmT0TPetG6wxrqz5tm/lu6fBmO8S29baJbN7rv+CTWPbk+l3
HoHdZu9lfKh1XqT9PdRaqKW6fL105LvKGub3IQZsMFy9DrmcvDCJSo6zXUgN6F/p
NOVJzFbQternfJCgPT1FGS99TR1Eqc04mIy+rcgGtud6iRNpf/GjL2221ImJvY+T
0bEkJasLymdmXNp3WTXfXcYVxw2QJizNZ77s3M38R1v+rVUXWphKx7uLcSMmiD87
F+7oILoBkmRZLfBvkr+zV3FuacMmHoQ7ocKMR0Tbwbnv4Ji61Gb0gco9X7gR1bH2
rJ2EaZtNnTsP2fYoPKW2czPTaUy2MukIs0kUorrsgAsdkYsZB6twkyJMgYGh3M+D
PeS+/hyLVOHtf378iLvi9aZIi/AcsY9Fdf3mn64ibiYIUw4FY3EvDjgDW3HRwn0S
jIgFWIX080gMANzDDrgvIOkHKZT2uGPBsO9qTiNtp+bHiKo9hYNZr34gCRTPYMEt
v1F5QZZuLO+PwfaZOWygsHPAAnGmCgOTyRtSIp8BSThypqCTO88kpYr1F020tiwg
C2mGOpWkWkmdE8AwNzFqRRDqnhOo0si27kUOBtV0BrtpytpEHmoap3CGDR8LuaVj
TSEuU0ZkR9n7PyzvSHWXvmGjHndWH63B+OslVWaQZjlnxH1Ub4u7I9P/t2WYBuqZ
uRINe1Vj5+xNePzyiUSwXLycROWPnIXXCheGBcPj3qx8GCoESsi8ncSYxVU7EwAY
h3/fayt99Ha+3K+5KKOdH6SrjTkcLTgTAppN5I1QZjNzgRc4P3XeHnZiF/R+H0k1
Ya9xRN9dh4TO7WWYl79rsVsSaHmg0Q11udVuPxEc68uT2ZBwDeyrQmrDBS3jv5tb
U88soNAu1QT22yV97KXSoLgx6U4lcbh5mrHZHVXGTJQmQzqEcEQPZ90ACXZWu4no
j47+4JNCRn7ZwXKd7n0PlgqT4URkKpV/3YDswhpbegTnv31Vk58NOmNq5I1Rk8oK
sPwdqszGpGyRtwN1y2nZf2q405dQHsPWgt8D0M4V2Y+k7HRc6npToBCvbRTbxICh
ql3DWafdAacBvAmxhCATOAqPRq9kHg4Zt/Gp/Pj9lGF5oxkw2WGlaGHJuHC1QTQU
9rE7/MOA4Grp2yqFiE9egiDX36K28Og9ckjLlPL0RVLTdM0vzWGUd1EbDoFclK2s
D3KRuFHNuiVSrQoePiUqEx/ikLdsE9Sphr9GynrGtOLJnXkdKWmUDOdEIjw/I+1k
Y+nwxcmJDKsY6QIVcWZ+9CDw4Ct1eu9HfmVG8oeN7QrltO4G/hpvbp+9Ytk26kSZ
/eDJT3V0uernnfTwPTpmyfpJqtfszPAyZa1oflvmB/m238llLGV4DOXyZI7W+0rI
Pc0uK8ws+Qu/0aMFKTl8VFA5T2CRabcRfZTCUULZkIIMIgVa59lNzm67k0oJpRLL
uOS7CUhwHdfkijdSdl9HVUNA788m5XsNg4JqnNrIaFr0Qha/342qyAecpwRBuKxd
amIlS2HO1urKHjqB+ESUrKQmhEfOaLbGzhVCKow2vNVVzgqKflZ3Yx6ryyO8fRFA
+KD3sb6L3QMo7ZdDOQ9Wav0SZwg6M7Mwj8v6fAL+nOcQrHtWe+MHeGEBGLgENKzZ
N2efrS4oPV8rSwlgjnqtgY16eC/WRnplS+0FENy9Ths9beTYgh0T7jN2bk/9em+z
EaAthegr4WWGCOBAcA5CnCbAsZvDvZMEsd/tU0ThDYPNtFn7CpgJrw+LnVFpMd3u
PypX4v4ZiUVWOPdy0z5MxO7JgZakdUM1fuxe4JI6Hi1B01VZ3h/qXHniUncvuEv7
KiPQY47ku30lrGKCm9C2+DxWGTLXmiUZM1zHttqwbKpMCfOnn4bDZ7e/pupo9aG8
PnKWcUduWYiTlf/WkXjEG4+BTF9yL6v7PWjDw5KlbLYbsq7MjNNGul4kY32F//aa
Ea0vN4iNPTgixY/dKi0J3kSXXAa35fnu8DCrtEcxB4f8xCniRfRof4MXVvPMBRY2
On4z0D2d2PIZGHwgYVgsYfaLWaI6X5nm9YCzele0aMGgNVu0PLb4f/+vZ6v8e2dg
R1e+uBD8u8VKRiv1xLsaasFspBjpawbNw5Fd6E3wa3GZlij6llWs/isWaOyWFjXc
v4nPiH95uNqn+ayMPu2i7ghlVfLRs05x6qBoAglZlWLQuCqfMYVlRKr86JJdvyaT
SVzL2tIb26UJChC+Ten/CVt91Dmiqsn8Fp0Wsh4/Jz1UiY7s4BUbYUIi+jVV4awD
66zxldnhYmTu1qvLKo9bbeE9mOyX7r3q1ebMsDs4FfqgBO7NC9oWwZqJURJbJBkj
UPUgb9ZoMtn3k5IQg0sQkNHmQcq7AKeKMZgCQjX0Pccm/YYHCZQGw1VD0edxGc9c
ZE6aR8jxKBO5MjC/7bDDh5ncUTk8EeoU33hOjkJ+5UpA+rBhA5VxqbmJDNxFI/7c
/HIJSmBTd5VR5qS6X9IqJ5qRjU4maL36Uic5IlDnj7Ze8S30w/HIjpLkwOqkh7lR
298tjTEtQZ/+F0Z8PQtgxJhFBAKimwiMndOKmGrG0R1ppy84+oyZUT5DsB+Fs4Qy
h1cuCxpvx0tVR5Uy1W+WUj6Uc/K/7lJmTPQLkYfjw6Nzy+STHj1Q9OBq2bzF8V4O
3qsfijuqahUYpr8mpVSvfVz9rKmyWNGvdLh0c5jPlkI=
`protect END_PROTECTED
