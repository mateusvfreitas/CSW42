`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
VYq0KXNDpw/vSqW1+DGeeTp+zVia0iadlzM3DhWKPTwg6WB06GhuHpUxslUv4VzG
+vSPjx9KuGWLsGFOZ0+rCMFFqRalK6pU2ykWoNw4KMt8I32+gL471vWF1N66k7To
2fp+CgUOxckoczO5/Yu8HGRLNN+rGYPU1kAScC5+LgmCDrPyyof5DOGkA6lIp2fq
ubuZ0CiUeVAh3fN+J4yxug3CCqzvdxUWQVXpSN9r8VXLEt44QYRnDoY1TUtNhUsW
93JULyjlZmZmdIZLixxribeE6xYw01hni9/gRdHwKI/pP1FZy6o0NFoquIny72dz
zt/MdRVN28gjZH463hf9eVHVbj7ll9Q4E+0wG0Kj0nr9pxz7iRDZVE0dfWn6lO+C
B++eIZ3jqKCdJqUErbzFSwJrMs4U2Z4k4IzkdiOhIFmS47B4jnVuWZ3EgMgIDEcY
Ip+1lCroUjg/afhyve1+IjQX8FfPXx1NNCwGsB1uJrnZ0+P5EUzA+Up/ZrL6o3mT
Ut5uCixyXn1xZlgqL5rB5VctqU+3aldCXJhib7XyrUCJj/NShGSzwS0HdAugO2TG
kT7zyiTFeNswac8BvPf9p0ll3kmMqg908BEfz3/hq/TP6hy7Zk4ckl7qFXK+lkkA
kLwtHko6cxDCrvEr0bSjcR/+aaheNLt6LTfL6BuVOHcClt2OWYYc2UTSDElWZsJ8
9aglumgm4xSG69misdWGoQOdKxqz6KgWJKN+fH8WTb6pQJAFp/7wVGHjNP2cPyuH
9ybsaPlEnQJJkPxC8y1cXZqbeqyDTIrWWpUQ+sobvfP0EYB+JeH0wWtpNxbp7atK
zPNTJ5ozNVI0W6XFV+ZEpBt5ojcCF+OsjSFsUjzacMYYp2OXGsemCoUrOR7GFQb7
ANwGERjIXD/ats9k/rayQ+XtLLd1C90LwlblA8JtEBtiMIOTJTtJfstDJjtePerI
WxgtmBkAmo9d/dXBiqf5q0zFr8MksuijXpeodbfcx1axSmX1jQSRWTkCsWlUZozt
N8p3tZ6/0Wf+esO+9bl2CJcm0yqGpdjgltFIPLgeGyJFjXov9qzA0lifB32ULWLS
cLUs6SUOEKeCFTMy7XO4X8BU2aWlIdGsUFNcqQVhbzBz3HuwrJkVS53Cto86SXW6
fUiJXfa3aADxZCsYWWjklYaKQXZpwwXqgKWNQbrGY/KD0gEuOYZrYzea3bsM6KK2
f58Arwx6uDBw+0GIklN3HbW9pxZgtru/N/znQdZAXU2or32kuo7NICDp6Ac7arMB
i5TeFu+astLmTUeXw6ZGzmp+iZaG1shnKY1e6Qwbv7es0t99GmYxiRV6tZqZuWY+
NQ4ArYF2G0QlPTKsbGvW7hVQr4ItAh1VuzbyJFQS/DIDpgTXq7JR/h9x+YVAEQiS
d3bhfaI7V1LPk0FWQIuSw3j1el78HTDGdn60q14pg+2BAMO7HYx0ZKOxnfc4rcTU
SIgbjwKVOnvlPoWnFyqhGWVVlvcUsh8+f/OXyQUost70JKai5W//eMa//nztb9Lb
cgB6THb2gGQq6/7uiapXqVBcfCQjt20YoLukcjp0p685sQXJI1hr/8uWjVJPfgLL
N6Eoo9AagionUlsMSdvGILbDR25hLP7DJ47v7Om6lC/ucMkeolFF3PWqiyuL0inO
LyhPOy4J5G8x9No68VQf3sRhfGIp9hsevGdP0rFcF6HjdBdzedrErAOU5R2C1op0
JHrq32ov1BafUEBDFidnJLLx/UKzxQgvwvM3f2CauSnJSs2ZnAElAHqXDnvqqdIS
VOhw4iENZPxRbwP7kXl7HnCO+KA46QjjrKQWLVWyCN8J5SEBvfAczStpmrXmiXDi
xhuLeOWO7Q4FOLwC3MIKVIA9nR6cxmyNthe6uXSLV9/4sz7Jc8qBjga6VgHOQ+6h
sz24MV04crkPPQ3ISpNvd2mzkgkkhHYrEkHIl8jiZKkd6Uf2IQdQIRLXK39pGoTw
ux00StSPZdIBMlPaPKtRKHzc62yZYzmKPSOxjMlivbV60kzPOrt86QUrKPlTJOuR
xBBpyQpNPLEJf/BsrrBL+4prenUNCAE+drQDpydDwIxWvwlu+68EaXEyKSxsJVqI
QpHFPbYgn/Miwl7W5ilBVousLwho39IfIl0achhlG7PDSj35uSGLbbkXKMS8XFEr
jbiaDWFJsAucYvSOwhu5d64zAHWCdfzHPps6fCPrbD0SMNs9SARBMFe4zdjACXuv
077FmXfwJ4Q6uHGFGs3Za9q8OgsDuSamI5p2ENK7CyyB+/tqvANXT1MIk3VBZNMs
Y5TQ5uSDCWX8bFU4VW8f5JGk8lOcO3rkSH24HMp6442yZA7OMuoElFBn0V360dfk
5CWk8JV8uyfjePo1vKntnOTEf+OhycV2ShMphCKyQQpiC1WMLyiOx48aSrXYHZOK
TbsSiUqSxXKV2zJK56YhnSpFJqqTNHrgnHGblucAfuh+yU/ADpxFySg4elyM1zkA
i4OL1RXLx9inPwgGK/2qlDH0c4xlUIhBi4oFZ6vkorFfUz3pJuGW09V8vLANiTZ7
Cng4QTFZiBphkdjeXQat+7inUq3H5f5aWbtG5z7CoIFa2/J4MfLKNvgVIkgdrWQP
TW3Z8zM5Od0Tcpy2DPNDD/5/G6ImxC6b515DhRCZfSd300rLhx+7+QqSQ2pk9qQW
Jdkjen6tu1h67oyOcBr+oE4rhZXaAmKygeinvAOpsO4Tt7XwYm5WZpqyktJSpWni
SG4mZHyPVTtQaGRON67nZI/w7aYoHzFfn1pgupcs1RG2UpScb5zbPXcxtxxJBUbs
Gx3xEKzzexGJVZpXSaIvPBHLaTRP6bHsKsKwSegSaL+ScGYdPv0oA0EFKOqnUilF
pPCMevkaQN5UgU+CQ7SHUEhDscwqGpjaS71cRH9HesSDT2rN1CTXAxJkzWYKXCZ/
LMrlqKzCSSfVyQn23jhYrXt4cixEcU9RD0hN/XpdSX2+BiZuGVB6Ss33JMY+xeJN
4s3GRwHWrBU9tdfRMT4ZZp5Tj5bXdwT6JB+Wbr0xefhOJxL6OZQOsL96etoPBMj2
32sywqSBzPpKTrpKoL6OzvCIVaCXMEd8hAPoqXn1Z88d/2ACLQOCMUC+QAJDTwXJ
c3ujqmi6rb1ku4hobfZHfVXgGoneryktFYRalwoYCsgcMRUK2C6ognA/OLwJOJFK
DplYILStZYNZD94X7hChWJUUcIFKimvHDZBwZrAvs3rt9aIzQO4pudMfSyjAAqu6
oZMQsjarQ53NWU+KZu5zoPTPg23pn6Fi7LZ7bf1kNfqarRkgnC8tpBQxYDXPGhPJ
N/zn5uUAil/N3U6qbkkWzby7gWnClab9A+CtZFl2JTpaNLMjmJVrkGTbjGPl14AW
znTqIql7lX2LASMzd8AcXlzS2ViuFGqnxcV8Nt6rWhPzAwlgNNyAsJPdjK7C6D8X
Uhkpenjdvm1yG/+98hIwtGZb8xSakWpE/BWYAcjh5VNlaegKmlS6MuurtOrOmdPd
b7dcBfF58bYU5nh5AMJJqWqB0E9jhNtp0XvEXGRsThKb+/A7rRz10NMWKdpPwbTp
5pgmI31IHzqzH9LpaQ/gcmmq+CR9NjmTBWNLxSM7zkR8SoVCWyp8qch33/wmlwTn
EyTvVL7cKw/oebYrkj6yO0PeZzxYEIZy27cB12B9VHNQN6Ydq9oxQ5h8OQqdWp6P
zx6kJtAEPTV9t1g7DFB5lHhh5EjHq8ExLghZJ3NsXzRFfr4kxagYa7rGfHdBppq7
CbJSOxG9+yiugxt4Ce10Upp332od3d61VshagCV6S5hz5PYm0SOG1OR3LbbEh6DV
TTP3AMpAofvqI6GRQhD1tjFt1LUsfY84KfPQ5X1Ba69nVb2AsYXyvoqFelHzAq0y
WWHSML7Lmkm3QkbuscLlY148z1Dle54rfktleFYpRTeknndH6ZzvMuPhoIWURSPS
nL8qSijS4dP0CA/mVFjrkRIkHZTXBlXuRF/XIMKq3j39DBgU252PNu2v41PCKfb2
71mZMwwA6eepoSmGGwvHBba4HQBtd/xREIV2IizbBJiTaBgJwmtvSacV6biNrXJy
oV5G496eXGzM+L/HN/omWFLg4QTerMw/yj5NqQBFLi6m2IrVW5nGfoQUCnqEdI58
qal15y3/xoZN5szGYNtYq9MRGbKJIKtUBg/rCgf/OAwO4CdtzmZGD+jKpT+UVawe
5IgmsMQsd+1o1CbW26TJ8wJiKaMof3KUwFuuP7DUlSRpfLxbMG706fvDfMov+e4M
VGAGy0MK1Eg02ieZv56agZxRVMtOkDx8lfKbZcBm5YyOGtagRwgLWR2tgr+5vJ7m
FEMZMKsREpNeuibG/tcL+RaSE5udNQXgi5lNqHtzA0rJsrLVDOm4UDytl7VIcH8N
NPDnQkImFFwxu3xOsZpaWBHUk4SSXvbDNSghX0XqELuEn9my2H1UPCc2L6hsn5fb
hQb5DN535cISzu8LvUjrPe/Vhqm3731fDn4kX9vc5pOjALE4/zXwfct5vONq80uF
yx8WhxJXuU9b6uYrIr7IPQeeLWw1TuDHdkeOSWTf4A327jZ1IDRERqyuQy9k/VFr
YX/4EmPqD6xT7IAEzPzCpXsea5aDqyHtNspA157IA9Tlewy+g8eoNTlQhJ8Sk9EV
VXvtI+7c7pHZn9sruDcIwXvULZt0/XiSk3Wiz1uvXcgS57XSSsl+sKXYnf9KPb25
s5XLa0sRwQ/o49YrtlkxXn5wIzipv/LFMbCDWmrW2ma6DK5fS7whB7WyO0k0ygsG
25le8mbfk6ra4HSY/z+OYZi1fke10d/ClN2tcPc7F/7QLn63avguoyzWvf/ayEG3
g0youuEBQ/3BiYx4JtnYpA1iuOGiBYug0mRQHD9XqbasYZZ7N4q2ADw2iasyLdE0
eq5HUz6UpQkdTwv9J1O3xhZPRbQ+nej/e0LJVe/vnMVLc7dLBP/h0u1tJN3p0J/D
KuLtuWPo66T+ZIdWbA82w6UxPZNcWvstBOr1D2EryfrMM75w7tnfT1R4kVIJST/C
5W5vu009IVPdrbbnYCL9CEPtG+5QEgj9QTW0OqyJekA9ARFXn0hguJvLKgzcWOyC
OtsIBanam0Z1szFH1Y4ka33aH2r0I/C5E9pgWV0R9DktnmrXc2ywShcts9OUlb7t
39BKX6wGOd+9Fsb6ZkPJaqfhwNmQ9kklAxmKZh9EN7grMpDQzDOV++1e74/Y1fwR
NaPk+Pq/mLGFnv1qdW1lYa8N55weAt4ScZAwB9YUjdXxxJu+A6B5U3nVQym5Hx2/
QcOFJkkhJP0/Cg0uWwGz/bDftxjkDRrNBWhlZn8Q6cp/IWkGhWE0NLrnOPNRTHpo
ickwzefiJa3++ezNzNAzoN5NG38MbyLt9tPfsQVn+G259u0r/QJNt32z1tMyWnHC
B2ZZuhuTRF69JKxfAPsIuZMur9lZr4+eoF1jqfRGF5EQ6BE8vn0PKpoNYN9tsM6V
Q8f5rOUbrdHlWfeIGBRyOhVKUZPiwZv2LJ8A30JrTaodAmPzkRvpIt0+jcwWRzis
h0qPq4MoboGiVOC1lPdvQnvl08Du6V6x1JvLxRdbfWPLv0hoROUtorCuFPaIe9Y8
1azIJ24wwtcZE54QqsFNhm5k7h6UIk+zbwzYJidDV9kaCGFTbdpIVsnjqg8cUKKn
WZiCDaHM3tePUpwU1JHlgdueZO6pmgXKbM4u6z6Oc6WVaI349nuR3ZQ5IUQlMYYM
ZGFjXxZvuRgpzMLF8RhIAZCNvqZDB+OVdU1s/MWhpyy0opc2cmR7vPyPR3RIE2G7
OaDgjXhyZlp/SqX1sYXT35FYbNtQq5epNhS1ZT/jpT9pxaxDjMVrf0BzCOMGjYZ0
o5rx46tM9AUbK+MOSNUGU2hcJtYsNXd47m1D46ImYBXUYqND5ZerYSToc4MZIrCy
iwhn6UaJrnqWTMHBMiaQYdL6jSIiuES63ZT5HK3Mk99uGnBMB3EHCi1wqW7EIO4w
kLFo7LOvH0FyhAXvHg2K+bRgTpgGZRKL33jOCOuAqadD4zNSC5JUTnDiRjlPzD/k
dyJiHHteahKtm1LYoiE6+3LRwAbk6JRmh7kCqvfjwR+AgX8JTM//tFN/+PBpAcVg
lwtHKv/hJZNigxD9wR9la9x2XV2DBwRyXMmIGxECw5aPjpZ9ibR1Bo/mjjxtmn/v
7I3EbDT3nkhFdlMiCsW7fPXvuSOG/603YAKD+TyQayE+fOaq5opcs/Nr5ewDjHFr
mLIKRv7vbW3G1sYHZ9hQdpii4BgpNnFom3jlz5h23G5zZHfYiPcEJfYT3gSCDkJI
mKfOoh0sJnhos2j8WaEvYFacRWy5/jBPIOA/R0Nq2kgZaxBOkeLYc/atXapNAIn5
mpoUJKQi0OxONTfIgre7LGmZ/NV/6Gaf0wM0R+HiXZC9piX8q/DUjzUHi1y0FJBW
n9i/K7N9/8qipvUw/a+wWFyVhTHjPZGLmAF5dun0fqpnfsuzzUomyM8NtYN68fA8
S/UZfCVMoM55IZbwsYsu/zK6w9BywXWmSdAdmRQjUD/aibTZ7otwzVxaInTTQNlm
0VwW2hkguMwRxzI9PZoJh7BK0JUTCaGIjkrl90afNaMTY0UgzdnjeGT3FVRvLu9b
mfZXw3LAzUoyY6EP7bi7w6KMWVEltpjkzqfPtN+LOXg=
`protect END_PROTECTED
