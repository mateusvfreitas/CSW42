`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WjPIOcSp/Z2dt1T1LatCXRX+t1i+VKfvYdmeUWJv5EFCIGVLQ5Kn9Pnebsrj7zPM
ZTTKY95a11GmHX6u5QWnTufrq1dWv8seOCazHMrMB9JCncdNywwURvFnUSzHucbj
6IkPNpbfM4UVbUoHho7JQITk1JjQRN1+jQ2pmptuagOMSYPO2I2W8bxGy02x18Vv
7Kb5PVc2yW6gP+hUpAzVms9nDoMSZhy1T96u9wM/zMGs1y6JCZz2Q7ePDzwxh1aG
4b58kmcve4zaveR81MMg4sy72SaJWXPzlWPjDoKloCq+boxkAGb0EOSr6Mysl2G7
wRYlornE23JXlgi2QUm8vJIyW1GyOLAUhC6Azeqgp8JX2rDVFp4suKOv36USt9r2
f25eGDt4wPTOA06032bLTPPOfw4o0WRvUYyhtSEjKMsbt9sUaP1E0PMvPY0ahEca
J+Xa67CIQeXD+tzh5gjMlc0T9J7lmqYUN33XnaPZxkCDpAMpROyQ7epsSFeo5Vrg
Q5G36/E7KzJBwwUbm+ZUDSlJTggMo0r//jt8PBcQjjY/oeZN7lPZ8vEP/Smue/Os
s1PdWXwz8vR9B7Voncqopl8CIjmTMpe12bUeJLGHaW2rP0PnN0QMbv1oVv1JUGFc
8Bdav9CsqjznGbexF87x4toU+GtmdhULJ6fR61fZumA9L4b/5M9ku+X6/bHD72kD
62+ST9yDCzVQwc+KCM0k7f2xFIdQF0bl/uuw56YKCELIoarfonCRkKEn3wrTlL4e
j9dvs2my1cqTrI/GKYAV9i8rDqpwCpzrX3PjUY1eMywoAp3uP8egDqTMu801zFyJ
RWdmHykqRWgbZRZZAYvCRRrWbnFVhdDzWOxoG3OA1eFc3MH4I6Vapy2IcxWbvLk1
56R9XysOhuzP2hRfTF8gkXnP7H8apzwNshzHGQ1aDIjuz34YLacIHbH/MgBSYRrW
Et8J2/tXdQxKfyYZY+YIsp6vhJVZ/m3gLQZGcXeLmtSiQb0YrwwQ8Ld6BGDnJ1TL
AoO915aV1tLB6vdQL4o9zZ2ZnZQJEct6N4LJTK5mnr/kav+DSWwdaL84Ll5QOMPu
4BAAeAoiYLlg/mmAW98jxoWtmFZKOnWeFpi3dxlSzUUwxhp0LbCkOcqUQ6wh+8Gz
VZkvpapYGebf3MGbbPe8sA772aDgDNIps16YUGad7oAynTz755XvDEzC1f99ptEA
SGUGZSwGDsJpg7VZZlI7/VEcUgtH4yVZ/k+30qiKcUfLG8GAkP1seKf9wLOY+o9M
9mnbnZtqf+uy3huOQthOWI4ad/DIJN64eHBSRO0AUOhB+XGr2P1AJv6ImCQBekcx
GKqnwOacFKMZ4xyRfATno1s3kGaejGFiOcY7ADlWDkmVsLwjpLB5IOwQWjEctYx+
+DaybgclcRNvd4P8r49PEyv8Blr4wQ9No4JemI6HcQoCmROitGpzQG1lgN6DCOCt
l5Mqg/nCSInzB//O1KBFGaMVZvuvKbsxsY+rsg3I42MtViPt4g09jmjwmwSy0NPy
9lc1zP6HpsQdY7XT7f3tX6sRgYx1WrmxZVKjVCLg0TroKak0136k7iaJutQ4uVuy
JylCZ1nOuSQghdwptQA43uffxy92m888NRIkmuZiPK1pMHWH8N1kmCOs9GnNtyzu
nYgl6ZO8ZFxGuENzaa4RMCQd2/h8WPqqAfodcD7OkjvwWRrK0wzzgGBgYFdJgDpr
LOT3h+qkHGEB+ixVSloVuSeMQE8xeJUE/RO7W3Jbr7JWNVfkmsZTKUzVbwK3VvTn
n3dM/wvhPpatezmzJ4F1WoZKFWtCY7/u41VKZG/Lfmpn7xuQ0J1KhIa4ygIHibnT
UHCkUyQA7arYik4jKoz7NoD/bpAZ8L8HfDl2HDCb2J6dGoYaaP/9vh0wxYIImAOd
aRKVVza7mhw2cER0xibjHlmmqtLt5hv5Fji1oeiYiJ2YaQWf+eds9ay4ISrAa7a8
0DAvqZ1UTpxTEw67ynYpnI51ib4eCqtwvIaEayr/jhSA6hEqlbFusPwRzHDCVA6h
`protect END_PROTECTED
