`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4TH3wkfdp8sgWzxtW+/i+OEdrlcUwHrsmxQ1JvFV+vFSdLsbZZ0gBuAhKkAZlCWy
dsxFAepcvMKnN7+VsaejJWW2xoyiIFndvghf0kvYoD3n0Y49Y16TmTPzVWdnGMGA
eg7BwnNJ7Tf9hA+JuOhPuR+zHDVtoQEAPB8vTtq013kBEJ13bUwQmazUdLMaAqym
GekZ3ZZ2U3UCU1ktFVf8X3UjZeRkbYmaYlwyeBPRZNogToG8ebciYVYmIcOdjjVA
x7PbXQEe/fGWviRmCdGJQWvcsfR++fVBgPrFbWm9AAUoBz6fJT4si7aTSu7y0zLe
Cssv/FQqBJDrcOahnhYTs+MLZHzgxIoZx+JxI9SquwONfXNe3xBBrx9frZGEPVoF
FhMNQBOm8GDIfkBjN9Fvz6EdQgfmvlOcT/pAFSh6Tq5Q8och12kO2w/YH1AwbKdw
72VEq53zYejC/Lew7PVWouChz5pgKomnLsoWmFo+3w6Cq5GTHXGiRXX6gWo+D6vx
5QQN2t2mDp2AG/fFNxBvsWtfP+2X3M/tVHI9RvbHy/0YCk+sfsKBPtOiDWkDPqoA
O8Bp7yJQ16ugCKdx/bhr6Q19xHerFkJoh24BUiIIz2zhZHx7Qm9fmEv0ZxYSQj6F
ywbg+uoE/wexqZ9ulFNS7OIZbGi6zBwVAABVeBKBc0MuC4aAFbCCRAqq/i7yXfQj
7ZumpPn56QnLLGB4wPOk9lz/URWK43kRISOBV4XRdmSMf7coKqhbduLalbryEK6w
pLoiTmlJJ97xGnzQMVT9CGZpsPWX9I+6ZPu3XzhZTRa510hE9/qPJatzGCopS5/I
THdpixH0bpX19sHgEKnGzQQtWrXd0gXwstVZatERpmhKqz1VtjOm+DUMHh2u1qHa
ffbztZKYr3lh+kgjefBSwMwPqaBNWHzloTk1FEEQa0q2yVW40B7Z1TBJOX7qCyz+
YaHv6BvvYtKYVKgUmRe7Sc2+DHd/S6A6Hn8VB87SAv7jfeZveO5WxaMUNgLRcNQY
g1I6AUhDYECN+KP8M5nqooA7rac8A5eepH+Qhwyzv8eRgxpH86S3jDPj7akvbWI8
MloKHrMye+Wth+0ex9oVomn8QVkWONGOo2WVKFhFGembH3yfxdsjIuwytZrbWiRH
Opyh3/ZVjupNgJ9x+Bm7XF+a6LM34malNaTr0eILqB3+ILNV3qbn66CVRnyNmie5
UGEkHfDkHRk5hNqP2ZuCYsoiyKDeb8GHQb8XbdUnUGX2sSDc2k66i+JruVmx970l
85r2AcCnGJPsEPD5dpieQ2aW7GX9ihIEmCRvIhGdOsoRGejJ6sPXxZqOkxoYh6Sy
1GuZ3NSETIw2+cvRaXrxfOR0lvGHLT6wzQ7U2mfnfS7mBfmMmYKnOfQmho4X/jxx
1JAPs/4e+L0z/RXIvVGMMjxtIr+VW/5zsPwSYpSFTkvisjCLgZXL1zy2zL9WlDDV
Ree6YDuYcoIUC2x65cdD6NLkrpx6B/tZihJ+n9y9D3XN207Afph1MuqYmJeGLlK4
LhJEg78zV9C3n/auQf1nl45aRreycHev2qk2vowJoW77jJ5Pf7kz3bTHtnQBPTdb
njSkUWFzR80S7UBc8YhkwZtd2+Wy95PMuV9Ig/G8mc5LsOKyF3ZCst1NauXE7Dnr
d57IkQ+xwjsnZuAsSLegYuswYPIx7pnoQVxRcvWk0cJZhmm5N1xXKceiqqSTh5nm
AArW9ykEw7M+MrrofU9Dd7P2Qu6PbkbPnpBI81gTSPlSWjyyH6+s+433lo58zSbh
DYZnX0vg6XdXHOjN5JKblcsLo18azy+onmi72Mm6nLtDKkMSfElWWf9ud/rKpott
MnV9U8cJ8jOJEg2yutyZH6c4Fwef59X8A/86+7wgS2Y44TTbPfcrkLcJMS/g6DEp
6EJCMACaEIqUH/KT0XDUdVFD41rgBfzGpnyzSSLtKAXhDzM3QIg6AxuekzCsbLGM
ayzAY8peZF43Fz9QvHt+LhIF5FPoOVcv9xn977rajhberT6dUa0wM3DJfiCsZPsu
b1RhhulD3qlXMpc2Mx0O2n4+Jgjnfc1d5fiEuxm/QydDxCCJVadCOrukwXOi4Kkk
uc3M92isnLvDPogLIztSBgcfrX70PlxN8JyYzC8sVC8Wki7uMMv0d4XRn1KfCAI/
hxBc+rLQrJJ574ChssCGjtbevb60kZJY+uWoMLppc11d/yrOobzs1CAHn0SrYsKr
91H1Hg+W/bz8BABtcvYgPw==
`protect END_PROTECTED
