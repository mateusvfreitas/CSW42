`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NCoQAW+vW56M4f7w1AxHQjmYUyg/UP9Yzdmlvpud4DKKFuT2MdvtiI/2Q7pMhFpN
rpY9EgNBW7Cq4hGBE429gZG29XoFCkaBnyUx16hLabAhGinA5bXuygYbXypuk09C
oJYrfbg2EdMAwA8jpTg6xNpNA94dHOaIPPtiuwXgGEaBD0G5/RnyXE02xVqGXdlY
KP3MQ5QmjVTMr3/h0pCBiSn3O0McL4WbmcrDN/JrWyv1fWBmjiRkTv6wPm/2pYt6
Na0F67l3XMb27gxY97gJa5RnHJJw+KL9j0g19NNpMn4EIcesVapAk97eX1+KrqXF
NRnVaHfWxNO7r+8+Q9JYVdc2mbyVI9gZFv0AKDpvRh0VKXsEMKcPFscpWhCXSb1o
Wtza4DcWp41Zw447mPxR2oNdaOeiTeI0pkehZoXaBoZVGa8XMHFKtC7XmiXbV10c
4rDiD+TAbLB/IEg0DJOHluQEAyhVN7/h2PxgjNaA7hZdE3h80GUf6M2vAIZtlPUN
3wW+WGUO2pW2VlIaYrPN3l/cT2niqurx6USu1EqVJSNK0koTIBtk2ioPp6bZbnBE
v+CZLrP4loSReZZvH8RrsUbJL3+zLJz80NZhTuoCX+vg+oELnUAcEMtcjcka84ZZ
S8dFn29Kw5HdRpke5i99QkJpR6GYbStJQ7OvUPHfw9o521AfiWV9PeYKHk1XMvjs
1U8davQXslLOeAGu5sxyJjAH4xUAGCIHhuRlMiarQCbkERxyRJPEgubN38X3PfIy
sdgp4zsCV8sCykAf+iVcV3/Pqij8inK0QuFTVNuHsM4osSYPya6WwRQ8L0XaJ4kp
O7+54tQs0A3fDhNKGzHObC2JwylhWlExgyINSPWSQGAHSMYEvYVz9JkwaK1hZhSN
ua7Q3SORFZCQje4OtubXl853XxQfNWhoDUCKm1nWL3/pa+qZp/76681ayeF2RPjm
cAz+I3WBL/2dTTUHx4GiPfnuSbXg6alopoTH4GnWQFoH1Pzc2rmL6sJo5dvXsAAl
ZTpR/Uz/csBwEdZMIcXL7xc4QivyyI5siA/B3tKLPXBcQTZErS9Jcmp/KAOn1YBa
CGqyFjI8iy+ayrWr/pLvcpwQF41YBZg2VI6D8YVpxW9fdUeBwowRvH7vg/LeAE4g
FvNf73WY7KrOuMJm8GMzj3LU/PH+Q3kDa0r75ViicAiy6AJaw2bauzW8frypRvzw
ioE9DnTWccsRNQ+7gbKzFMAqnLyKC0IoKDSseOxkCgEjEuQrYGNI9AzORh1X5Pxi
Qh2jEHFrFKtVVhwqKaWk28O+fIqMgydrGQmLpzYmQK/r6VBAT72yaxfS9hQJeRLr
WnniQUOGt0BQ739vM96d/N6vblSWc6BjbNjzN+gHqCrdwgoEYvn6gkKvlCu6aiDA
bl4eh6U5sQb7I2hb1AZm21lHMfATZn/f1lTl7QuQFVnbsimdbDu8LB53TjNuYkqH
lSbAOh4xHwsLhWymSqu1cZOJUH98NI/yDdjvjJhhwXz+hL7Sid7adCjOL6W5hqqg
we3MTlHZh9zysFWeIgwuNfQY+j18HNqD493XwgQPEwq4ynIos5sqBenwRNW4mX4G
97ubtkq8ovkztcVmLpOhycjUpCG/W1uio9Z2ZTmaA0Pmsyd9MRX08zurjl/1mTvS
GB9TLIeHjguIodfzlRmBMnmPcxYg+ynC+2FZxU4TrA9lRQwaEscR1z7f1pAGDNTa
sfJf3Hhd3OvaVOFxbuFfwtgMIBlOyRqAuGNgxAg8y763ExrEryCKFLb0G04aH+Ii
K8qUxHj0/4CwMUnz+h+9i7hGklVsXWadaPpKl3wS890NWN6iXTVhKSCCiO9cjMwI
ksdbkdbIeocK+0pBvfklSxUeB3X4Yp2x+e78wjMZDG0CxGF2kg9wjoquxzjjDU/V
y1Rzqdpt/jM6r95K8tzsNyv1SN6qnqh0o+ADsHOiYBEi8X7bjiElncJj2Uzkobhi
qi033jGS+iqKLvXTRgpyzEUpCG+7EfZLiVKoTqyhCTsUEYHdVwvwddZaRZlpgsZr
/X8XR6uaKNvdultEWgEgbKTIY86R0yeHNRnpRXk4JMkfykm6WjN+irnRqjKOWo27
6nj8HcEXS0xLL6sZHd7vwteT9IyAM+ciqN2pBNkkZaqFLGGr5k2qa7timIakiGtz
QL1f8RengRPHeqbonQuDYrilEn4EHCNY0tchn1YIxlQIBJ1fOWeDbnECk+O89/z8
BaQ1WX7Rq3/iBCsnOAK7GkbovtRYmB5sAduqIkqJyPdNT90Orbx+F5nVkxJdbslb
0jV2B4Xq1/5PCCAIxXRpYxX9oUJsWQNktc1J26QoPXY5agBzE7CjfzJrRxhaZe6E
CsePrmBExHASjIBw+GP/bdmQ1otZiHPxiGeTQMPFrpf85NON/SJmEtmBgkOQXRRB
evrliHRZh6R0C5FQOJD92hxNBao/MprQ07cwbngFojn2KKSGnSCIL+1rwe6qWN7K
U7xMsbAsBI6DmaxW1suIIZiDDw7twxyokr5loNoaUH+ESq826Pp6Z54ukwXPx8Y7
RkaNv+oEzZbN464ietdCikRR2lDlqQMwODXn7Y5XNDcskCINjxr2kQcDvViDTQ7m
RUH+Bz3syhBnCZa84zQREpUekWleMQhP2wvFn4Qzo+ItsRgegv+Rb1XnVXbkz8CP
hSKRx3mxumH12jTmaP2at/s32hiQlPlpc0eWE0p6qbeUSbLUB/GcLnDvD1jFrABs
L5ZTtr/HstzHSloi8lbvXFHJToGTj564oe7F0YB7WjR3keN57FrUvwDixIOebOrV
yyTMHbMwTOUStWKx9T8tA4uQJpfSuJgHiLMgYGat9/IjgFMeNHWaTFIjTvYejV49
XUXpFbj1hSeZ66FxGSsKM2Rc/0/aqxlQ+Gw5gKx9iQzK0izaxbSFc8NCeaMZaBXG
IAbT4eXvT+BZm+5DGfafeRuJNeqrGekSRGs43/kORFgwpAcxmR7cbBK62p7TVxNV
UE5zzVeH/5jFxfsU+MuFA91Sz7YOZYT94NCAw2Z2nftBCRXiwq7UmWmJ6DA1P1Gt
A87luCt923zTvsI+Z2j7bx+9SCfGR2VCjCLS9YCMz0sdWa9W68Kgf6ySfXI/ooWi
8xVXBCHMeDEpBRTdjrTjlyddfauotHVGZNQ1bKivA1w0RkhvNmtLA38TCReRVpWa
TC3h+k3o/tY73993nBWFg3Kk1H3s5STOd7yDbM8Vi885nnX9fPilcUE+1DHniU6A
+CS1ANY8+C7XJksPwRk0QhsUmb89OU5kkIPs5ME9DurNj1qWYoaIXBjOUjOnYcvl
qDy1PKJ6nsHxQ0HHGU4uD4drTkrI8NRxyYDVxXZfJtYUZFAoQkTMnGnqOqL52QBF
yNSUKDpTaqbbl6qoqsaTgp4qL2005yNF1bP/g0B4cUVPVUGDB7J/1/pyPlHP0GL3
9W/lYDBBiGj1Uaw8iYKvhvOrZM3sQQqvSxNJl0RNkLihkiXccZgCxux8zaoGVIev
dHN/xCoJyjoomM0KkJ9/AhYFAarCDATUmF2L+iV9Sziq0HA8Y/NdZCInXL/nlPcJ
Be+PMxdcBCYQPneF7MNhVKPPBRJkP43uVEvhIpL2EmAwDStY/m9EXXGVuGxInVaf
xCoLcUWV7Zqgl6VO05qf8q0ADw272MAJWV3IpzLHwnerb5q3/VbPJJ8dkpKyCmz5
jwbjpNenFkl1CuwqbF1jynlDoBNEstWRfin8kCSK5AjWArNdcczkr4E0ksM0o4zw
5ogLaT72EdNp5r4ddigeAlJrnkPSiGJq3yF4YAWuHOeRePuT0jxPrCD+ot8+hPiC
hWSE7hnUBJLNMavm0WJmgqyHFX6q2gMrUWWJRrM+aSRNZTDtVjUomapwYIq9nc0C
vz6MEMh7T7FdAyRrCQeH9TCad0A/VvaX+2s0qbuW86RtBunvgkcKD1ijhYjNIdxH
RfUDurGmhsXzmrR6vZS0S1d27oY9pNXl5j1CnCXQH63U/agiTDFGt7VcN1tkKiOJ
xTFcXGyZ/OSvuaqfbccmH4SDAmM8JTnuZnG8HKSQz3W0nq0xpJttit0ITRLFAz8Z
vKm+9lUnJkHMJN51gacIu7Fk5NMzMIf6qonw1+93AHOmHoXjH1Ya+5mWfLagjvVi
MOyATCBX8PhSjTXlI3mXYHLsVabON/3QvVfZnoRGPQYpoyRqpcX3Nr2PMsAvE8jW
CNQk4OdDrNmYx/oRrESeQKPy/0RTkJ18bfHfxwPJiRQd2TKkm/1pVN9nB/3LEQGN
/EPMaxfg3TfxBGDHCIHKv7LpBhNNyejQHmB7yF+HJR9VnO2cUDYVs8Uct5Km0e7O
aUjQQrBPh6xWNRXnXs4gegDj4Cvm88BCDoN0sccjYdvo6gvvQysh+oDG2rpFv/Wm
CvUh0Wj0BVhwj5+zFQ3rkMSlC8bYHGyST5DPkKES+kmW0KMWUpAvJJWLbYpC/5a3
oioN1MGMNBgtRJz8nygc8BrvjQXzS9jDEdVDvLIrTXFXzRM4T7Sje7FXMbmzkrAg
99o+GDNvxkH49c6CEy05GsXYb3oUVI4UTzBztvkiOpp3pkcdPbUJnRRt6lGCXsKM
rKI+aDta9RDGdeIYqTRSZiplJZ5lkgYlEu9HzxD8t8XhamJw9ibdeCiKliN0KyrH
sjRyNDhNUcvBp5MJafgTEzhA8oux080htnBaEh7l27Vnu2ni3DjZP1o9L2g7yuA1
tzxcTmcyvxr7P7TrCmxtCzKotkGAvXT7piVvxbwuG6F2+/YPQBvhaPNJhkdxtgGg
T8M13axsvGcX2KFnpXKqUVA8LDS6En9HmoF+BHbEaTxyYqemnvt39IJickd2TlBX
kbFy6iWfT7pCmUJjpHPuqQ5d2Zlxdrh0HR+WpzSwv/TsnMF4BpF3Eflky7GT0HtD
CgZBmmR1uSVtWCiXGd248E2lezV+dmQGBKLExxgI3Nz2kOxHzM/gr+7by4N9h+J+
3y3aJN3/XZ6+W1h4jfIvajDQExL1rfjV95MZSVmagNQDq8occZZBuOSx8G1iJF56
acWSaB1xypPx2h/EwWgj52fDhXWQGygOvvH9BpowWvJjRBUi/Ruu+ewS+H0o+DW4
LCAIFT4PzfJZa7/JQv9U7EGeSeaH2YokpcCzWfNO88FlLoy6CupYb0+iz7eR2Udc
4zyu5JMPQMZQpe7W0XPBYW4pNx/ElTq3OIq9Yo/jI5uTe72CT6PoKn5AJcuKPER9
HKLIAX1Q6jnu/cq6sWafVGF3z+Ow38HCun4qmC0vBjD8LyBodvoAwiRwWrLTw+Eh
CiKbdUmrCpVHORZYJMlcFzaMJYljjsswD/yNgYqvN6O6cBuMXND+Rwm5/iKl0lY2
uSAqGQA+ZonV3wudVc9pURox7kIZN2Ousls6cqo1LSng5kg3LhIcbZEG1e0HjXSR
A73DgIAygWYvoZxc2tTT+qROayc3VMBY5WjuzIRh2qqxiPO3Y4PZOQJE5G/JTfov
ts9HQM/5rEk2E7VWw2Ks5gslcRNJTuYCdol2kTD6v/QiHBnh3t0S9y3meB4zNBrK
FRZgIFwj0jGq8IYxweiEjLLhr5xfkKXmfwzso0XeeaSUBQIbHjQ4ctcoodU/1y8d
jD0ZafRuTcGbuIICSHcCzu8JceCuwzc7uLT4s7+eOD9nunXQlYHCGpisZMw7xQEC
Et++pJwVNSraQ40otrfZd8wmWqBDT13C3JbpBxyogsfcLr//FUATchK7IgRIhJWY
iRCYPYIvnl4HWZNRYaqF/7lqLXhCaDKCRa8ILpY4KVCTb0VyKkIhCdMU3c+t9VJ3
fWU0aALjHU5zQShDofiutf6JQtvveFrzx33EAgYYFtiED3KGCWVqdugxSAsI1qsx
QSrqzNcMQ7+X1k/PW4E0depQGiOrlVpQB4yKWj4pieedM8Gn7oQ0vcWSlUyoC4c8
cOBKlME4dAjmzhi4hj2vb5lPvLD1aq1MEnivpOE+zLwkZwCfSJrg7Do0bSkl8LrZ
/mblLJ8SsX7hjwJsub4gXcBOprrZdl5Y0EFwImxbyM0=
`protect END_PROTECTED
