`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ApeV87aF4G87cIM/45DjTwV3DDf+wMIGNGuS5fE5/T2widwQAJV4lFIRz8I8VdwN
pxbutzdLOBI4MD3n4EOla3xmUEJCfXIT+mRwB2CsrfI+xPo0ElAWzNq0sMrcvYDk
Q4us05ELzomMyZhSg5qdh6u2zBiCgGMDXqpsE+iTE8ll5imlmApbZ8+vJamiS4Do
+CCap/Hu+cIPGmX+iQ+m6KH0LnFLe4dzENTNTACoWO2zeNlwXU3InA0w1CzPCYF+
jzv/Jj0p00HBYpCVlKA1mFD3ctz9u0xF21uYhpbIF2k1ETfi3Q+vPIX5vvj5Q/kl
/JzprGCS1ibG9UQ/mYlV32v78vlvJbT70P8fkuwSndle8mzAWWOXwfAQ0/i9eRCa
RVMVQBSyu53eWHKKpzbEnBOT0/Dz6i8VG5CLErCUxWVmnw6gURQkOGva7CDOLuaM
iJt3388XNVpvSvg2gUccojLsgw3dU9yYKhn9SKIXgf3KUdkTfMNnwl6/Jx516S3p
l5Uh+ea6VPRatBTxIehWnmZSuVSGT6jEZGD8tkEildUhdfEGMErxivTm3fPer3My
YoybT5Qnfyg4JOX2jYmr8aac880NsnO9WgCs368hkatCTqdZAYjBEH4Xu5M7evo7
fdEOnYTMqnZ88XtQ1hAW5wKdK55nwXIqOadp/MCKSHx8TPgy9kTnknww4VfbBBNt
aQJP2ZV6ytUBSF6hybe6cXrJixRJH9Z2ZNIEFUkoe8NfFIdPbI2WuTW2qrefH8MX
kdaIKyiXzyPjr4P1DDBjhsofzfk4UWfJI4BHCCIiOIEMI8BzRpEiu/L0RJXobJpm
EyB9XAJyIGWQbKXbqDR7bPrM5Fff37oHEd0I6nrDjuVcHHrFVuYX/DUk01c1MWQj
HsCkZT39Zah0Ms8wdo9toW7eEC6B0W4dN+awpM2ABQXrpj1v2TwUeD3FlI+8Ogza
L6ZKiUhWKOFKVwkl/4C9UAQrrBgU9GHyDglKUidXdajOQm0t9OWVhZmuuwm/L9Un
D3PAddSpyLRcmB/4N/vh5hOVKBRryuXQh9DqfD+FipFLAW7kLZPYx+S7FDVNUqgr
A4sy+35UOL9+rT7hn1iHM/s46gMhi87t87N5cjGrQfJCjxSYO1I+/0o39xexI72I
TF0V70W8wZjESukwPyeyHsSNVzIFDmLBqpAscuGwibJPIM6Uzg93gwtK+5IZKqxA
3dketrcYvb0gXjYZT1UxXgTVUD2ss12UDHo+qtDOdJPzJe4gNCvyOfYQCSMihAcl
2SYxhUKxjDuL9RDm+zbG+y6qm0B3cNEivxI5d8BRMKgQY7RL0/fF72zXuvJeOGHC
Spv+OJp5C716lmFgdeGZGcdqDsRuRIHetK6oz7pR0RhvG8YqgB2eg8KVT49XUq4c
1lzf+EtoHseBKHxhkSpUPrVh+NURCPLMgcvYbBOXN6uPfxoh0eLx3vGa5QEqaUTr
Zji8SZASLCfMGXfUgru+yrJgKFtCFHw+m52O9ExUQcH6M1CzsZ//v42CiVtDmte4
1ZZ9Q7DJPANjYMQc3CHMsV46UrV4FYEw3fWraLA2xa5zs5gtwKdcE03oDv4NTJJb
CajkBRWH3CqTXLA+nyAZsb9KT6+N3DX8Hg13QnvZWLFUdZum3GpCnpcEzzUi8Ajv
qAwP9IeS9qyTnkvwrw73FwSq2jAq+cx2tN3Vasg/qCjP7zDTS0wQKTyzLEjxeigT
IWhMvUXV8lnag+StugNW9Hgt2RqI8JaLFUdc5jKGKdT0pMPCGzToOD6bRXmuVnQg
CCMxNZlK0NaU9IVxObXFJIWaMY9lDFH4YHBNJPw7Jk6pa9J7nWbMYi2GKzPUL8Uz
m5SzN9vW5tbfXVg4tJ9TomZlIduZkNfsPdNi1Cx4j3/n9ajkWaoFNCs7nJo8ZTSG
ueiEn/VsCteGxrNH3NH8gH+WKyQxLS6nfFA5/UvPpsijyEtmCLjSuVjitnVE/z6B
t+MWFCxOJxouHg+Y3wihqN1yWDqWbMEegv5d6G3FDrtPH9hAnpAS5ud9mTlGMefm
Pi/5xf5uH/O2AFwatA8hHlox2o0BL2eI8srJJVVEsEX9sJGkfQkO8P5g9+je+nU3
nS5XITriyN9M6a66YJK6cN1W/2I5gN7t3mjraQ2EYYigXcPdekurQUzPeSUyvUMM
IQHMx2eg5SIR3zRYL1+OMZ/ldgBAcHd3Lvm/mO5mIJX/goazF3iS26sJZCsMcfHE
zuzhZCTz7TYIeq9uW/7GdQ==
`protect END_PROTECTED
