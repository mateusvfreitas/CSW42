`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bslB1PXW8k4dj7MNNXiyoOaW+FrCOmnU/D/RQIu55G1rkyoUqPQivJl1KKGKdH34
O9PMcR+xIusb0uUaoLZGpLwwhw7aJHwmbpfRhwm7ETfppxOW/UgonhpgDe1+7RUp
zypyDICjt2egkxDTIHqz6PR6N1ZJY9gN+N7rWSYhxjM9MEKMbIThJZ3DKQEufMLc
Jcdrb0QKQ774448yvf7jny92YH/g10WJTvO8auceeCtVn6EitvbIjbdEhXb0C/5o
EtPnQHcZtxI3CHNk3cnneLW7eKJy5KwS47/xfA1UZ6N19bBW/+UPFUENN9Z3bZX9
kZTer1DpiA7Fb8CyhAMmjymVNKZqJg4764e3Zr360CIE8yg/Gj+ih/8yjZL7Qcry
5mjHKMlPa71vuuFDgmHvQN6eJQDVVeq9DE09BroWFrXcSuRUlGU9NDFSWygYqrGu
TuYygXWol5+LWr2ybSasSjfyMHropWHjhBTGBWzLsVVZYSxtYeHlJeuVry433TYy
QDsxDoQ2qcuzneZzXl59x3KFHVIn/qh7oXdXNkIfwxmPBMoyo4xyNzej2DVemiHI
4mhO1ib0BOznqBYbsIBK4za8xSXjW2PwgXusvOHTdxPPxqg0MMQXa6tIrGTDs9Js
qcj7cm9s2ZmFZpgpURbwLaubQVfjWQNVPKtORQWBoTKXJ/MtF4aSQPY4rzvSifQG
zPuJ60a3J5qo7X466J3thidTKTAvm6STomHlNOAq+3u0QVNoWZNYHlx8fcBjAwdl
qbTj7xswvHmRAokGDVDEH9Jy9RqDjOTVqqzPQC2oeJKqWdmY5cFaFhqp+TpcvjUu
n/pkRg7rnS9pyqxnqTkkelF7Y9xvDiTMYAXPSmaUTm4iczdpC8jO8JMFwmuULJb9
tqybu4R9Y+LtH5lRrZByB21IlEz+8gwml+xFXOfgujbbsZUi8trRbUzskRzs6E/2
MHVibuGx4zFMbsxs/2A8/3NqqAKvR0vBZZxiwhfF2SLaOROXQkd9r/YRxwBrzM2w
8uQNb6OFv/w59HYKrBGvKOi/dcTQNvARiiOkSDZbinSRr4kLhO1PvCPJAB4cgC9i
rG/0dqHQeYk7x1Breax+T8Ctx2KP9p5UPPAknZEeHEXRce8VQYUiSbx9AIBlwO7V
hwszD3uYzF3UUOeTC9uoELnzMR9+FV4AeB1OboCOwLqW/rihdIb7wSzSzwk5Zk/l
Ym3NRdrsJ+Qdjd51hO7Xvy+gMOhg+FaaJmuaBVpoMuUt9igZKpsK15+9eoBwVPNW
FqK3PJWgbzrsbqIBwHtZPstQvH6u+nv/aWA3CZZrOdQNFjxbJ3CPqwgPlytSAPLb
PZ1iqL5IhnEAU2avGSTn5vkuA/KcttW9S6Iog3v5Jw2Oc0GPjL3vUzqelgx4A7bo
xpCZrru/lLmn+tIw5x46AwfLcVQP1s+cN07OZuHl0BlDQCR1FQNFe+Iz1s21k96C
5aTRq52oVlVKeBHnFREjX+lk9WB/Jsn0t+CwVfKAR/NSP62jQBu4dOVvzZH9Mzav
7w6DmldoAuMlyaaeeOO7Cue0r5ZEVmMXkU0bpg0d9BJz6JndwMs1AbLTuKsv8QXI
XNFMNJHQ1QVCzuekqz5BaV+1oLnEveFDiPfmJ0jramAWjCopRReE5/7bTg4IToW7
BvSmQIe71YYF/iHdkXi50m5+91s4UmNvTgftZ17iPlmN8D1g31g4EAAgR545aRGZ
GW5G6uQ8sJvNmmYQAE18vzQu+7cYda/Dj2CZn4r67PbGD3NBGEfzvT7/XRzwGs6w
mosmuAYvgr64EOMo5zxWnedPrtWxaBO07vrcoa0seZRI4hy8mkAvWtsrxJWrf6Ds
xBCIpkGHvwtTivIChL54UfeCVF0KsOuLVJy1CLofs3EgLhA1S9ZjrNDTeh+Fsq+w
XFaaDUpz6sPhnN7Am9WsdLZ+Nx6gHLHTF4MbqX7caqAsaeqlA0qg6y0SWHHrZyvY
0Oly2WJd6fV6aDVTomIWSYRNXAnseP1jm0Q49bbTRb/EwiPucgC0Rfpz/BPk4k73
arkVkvaVbUZeLiBJS4vpyjvV8JoPxeHXslurADDVjLJvZlU3v/l6RdPm1hrtelo1
zMb6XxRWncf//Z+YN71+iJnbEgW+KWaSpuVHpxWKXcpCkEi18XOz/G9NBdzxeKyg
0bT9JU9B8GGqj/RsIEraDoNJAVZdvQcQrpDZKlWpR0+LT+rA2aw94MMlP3xTULDv
H1bj32lGdBqaDF6XAuaSAKAaySQL24xJo2rIegCLBGNcw+F6ibn4PON/n2n8SzYY
n2ghSBHQmc+JZk0eKFRu82p6XyPdcMBNExBA+46CQaDiSBssamyY5g2kjRwBRU/N
ykn3XIz5/TIVa/aEQ8kQinwfwBsNrBsbA/nWcZxV+3/TaDOu3ibrxaHSv1iELCMq
/hukYrdrRgPjkZEhAnesOVut5+MiOJV5txmq+76cEQv8rZ9Q7XPFkLODIlZ9X7sU
mVT6iLnpjN9CUbSLEt+MFtmFbPALWnHkyXP73YWuGvKWnRwbUG9OVjSzQraeB+yC
Qs3O4utr4LPTVdRKeAOOK8uB+AVjIlLP8Vad+PwpQw0tEAGUnwHzCocqeJAjEbG2
1awgiM3PLGmIo8l3rTsh3p5vaAc5bLFNJ9/K0F8EEywlyZaE3HIkcV+d8l493Gqx
y+MhO2fReRv7JoQh0K+MjLBgyRf1MDwnJVzOBwNA+XjNYKFccw2ZtstdsTwCOSEk
2R+NbzmEj4reiqu0nu7Z70Uijx1AFcgIcjJ/xUlNoleiJW2ihbcNuCEnYBwW/8Aj
hrjtbpVGKugjzp1K3xu0OFCusVW7fU32Pb2lBZsxg1+PCqRBuk41oeJVaqB5AuPZ
bk93K9OSZc4p+o5I07HMchrDIB14iygY3ukbgssJ0q17TwbJ1mceK7cNpYEk8TMH
3B67wb1ngG1qcR1+gyPQk2uuA/ENpVD1VONEPUK2j783XZ4Q8h78gJn7Dnte3I6y
is5MBCxOCH4GNohEfEk/hC96NAXJZXB+lFdY/RlobajrGrMamogrtcw3byfZoOO+
r4js49DcSvjKxvpNKmYhIB7HSLYo0syhmOloyi2uZG9L2YtCehJgW+BGSxg8Msuc
UmmSr0g3x2t7UQZ463dOIvvcA4a4G9QGIWu4YUZqRZPrOb5NM8kN92cYP6l0DJV3
YkGK43NYrpXlLy+wv7180my4b6SoDNjflSPvp+qjsGGGBBpB/VnHQRVsMt81RBQ0
nHim2OjRZPjndFaX0q3k0saKTp9YD7S8rwLydamdtwbBalePdJHadLDeP+aACcad
PXMhT18k3q0K+7oQXCQ08Te6PIOTlagt4JjzkFFo7BVFuc+teNBgMrAum9GOOmeP
2DkDnvKTIOjfVNuE0mTzco5AJGFH9dOi+HJOASdU/chcyE/ivHgotRhQ/W8Vqm5E
mV+38BtNClSQqk2drOfZYPHMELB2RsPOTykMUgLp8E0Z/o3noCiuWXbQDaZ8GUhS
oZ8H2t1ZhC9K00PWtN4fnF/suM5jSnpV5HdMcyvmC4Pa34ZMUa6jXpKsof8DMPrt
Mq8qBwjYaLgXjzAujCfWzLtga7nqTF1Ef89/H87YaIVSA0cq/PnhlAWDZOWj3nLr
udqW7aUWuPnhIXU83rt7UHuUrKCWepHOfuW3AfwDP9sUmOeTmqPY4/LX8D9qrusW
E24UpjuI6uPvVwChgZRZR0SsbFcpmXkz/10nEQTjFvHmEH0QRPAm/k4sRbuqYPNw
VpHsoqyHsbxF53VMOky9twtGidbKduV7EMWxwpmYE5ShB7mZsW4cUfX7V88auDCg
svJ5oMSG/HGE3uMyQhYUL7MCN9tTWcX+LPwowc7v5BjDHR9JMb5tyXNdT37zYCy9
BmiX3jyUlcrNojNFlEs5F5f10kFK1zTasqHw6TIzuT/T/srC/1Km7CY7PlpiGDWM
JCCilKR+SANiJMqE9rF8xDf9xeeRGFX6aRt66O0tVwgDMkI3ZSRCML5HvGamPgTW
Bb2rRXX9CYw8mRrL89yLPgOPLbbhu74SZW61jCBkq6w8EfraDyp0mjr9DgEhGLuX
CVQrSS3EL5oPzcQ8D/MnRjM1a/d7nPsZJCq03C9fr1ER6EgjDg3SDBbqbVDak8Xi
DNq4XD1j6yoQmvnEoLgQaUhtEEMZUjrwPHGd603HY1kVvsanZBl7WvJcYzlplFUL
FeIfQOvEJw2FORbBvGt3LpKmPy6phoPJt7kmt59mYc/1F6rWxaK0TjoI/guuzktX
UiUNLwhreiLBvNctRXg6coV+k2Y6sAhT2OV0ELsIlnmrE0C+/ualvxkk2NoVIu6b
Ek7jq3qpPoxgRBLp/yOWrN+4TD3x0Q4Sb8he8rD2fTgQVYb+5V/SQnm5+2DzF/DI
kBsXmRDi2P7MuQ//4SUvHp1quBXIRixyX9HLgGUU/SPi3y5VWnxS5ZsAld2LPAcd
8LtFdVWBY9s2+UYoRO48HiI7ahLL2/Uck7dNcQ57ji5MM3StzkEsXZoCWyiuaMUZ
o0xnkKNGXLCZKDzuiDx3+iPqwogNB1jtN7o0ZA7Hw1Qv9+T+m3h9H6W9oBy0W3z9
uYS/mGk5sBM9fkOeQcra6HPf4UD4yuaR8tWo+zzqRZrfOwEi/6hWTx7PH4v0BpNr
ejtKGWgpj/UgCQ3chVKCWLYeptHwzzmPUGAt8nY/8qAA1PO0bXLCRa8fSK5xo/Jb
Fy/nlQ5DoEoP2anI9ohgf5gu3w6+azunFUcbkgNlP+R1Dqhth5yuhgb7/pV33PRe
zDcctvLSI4XJMwj5aNGJv400Gb5GGDmMs1lBBijr5aLJxNE621SNGR6OGFmmYdY6
E+x2Pk4i8jHxkNr6lWYHpRsk563483P/BGefG7ulTK26F6q6ZJNIYfWTCeFj8RtT
iTvivkx0y5SnKqcBq9R7feBf2O0ZBbar5y9m3nWm9YsFb4Rws8AOcvQ/0AT6FBY2
otxbnq2g1Di8LKlnqjJO0Tt/1DesgP6N8bdtaBELt/Jy/S1dDCmuFdHQU60WhAes
leesynGcvvKiKnQ/iww6okwh1OALCcUh8PSO39SNfZof5UTfR92oiIsydo8xU/tG
W5qRyYn1K99N+L4ARBj+zbcL8yd3yFNEEc+Ma7bWPlA6nWjWOl2NMwU2FI48VAIZ
WzD4n2SLeSkCp8WbH5lBMvT47zrWaUg7Ie+muJT2oEkvek2OJWQspNfSi1dXUCBT
v/9Isva/+ZUYMI8CNirk+gy5NGqSnGZ00qw9s0xHzK4gdjTmVsceUjABJDw2Szxs
yO8C+YqI377vU1ZCIdMW2FgoDqbNwc6u1SBAm+NLfU8xVNnQqInefgCdH4UQAkkC
60kSGUZNP6HMRSSRyNSNq/OYyHUMPeqMfazkmgEAW2UZ4ISD3HowG4Yh/lQKJYvo
qv/2Mm+xcrguaLfjKMZvKSwVjZ2xXFROtN4V4qzQlRi+hW8DFIXOeGl6JsE2RlBS
THHrUkbz6u/B+7RvigmNEM2XXjSYyEJK7y9D0azhPj3p5H+ZAN9g/4R/gD0qefNh
KgeZ7hh71d8lFZI3KaG1NkLIO8xjk0AZ8ekNSAcCOlglhCHKfwZEZugvDVmUcy9U
Fb6Mps8TcyiDmdj4gDmOob7/A+4pnNbsnusOUgrk6/iS+1j2ApKcdabTNauuHVQy
U8E3diSmLO3ZAPcmrMfs86QBjzbX+X0mTjjZ2lt660DCN19UtpNEjG6cUdFPkHHF
dwW4QkAFyK4krSshkqwmdGI3kH9P5fHJsitoullV7grRVp1n1vHYuCyNXTgls9k7
jDmr/a9SeZGYAwbNB78JixgYCMapPz4HzUFoh79yuQVom6e15sbGapJmpSN8q8cd
/Silm/+UN6rkrvI6MByDQq9q/AQKk386th3u2lyJVx2t+3j1mMekFoxznRoHkRsO
03j2yRLGA6YLbi9hHdiFMRkR72S4UBUVQxrTzgNO8ZqSJ6MXb8yYhZ+OvhtkycmV
suNSlgvdPwKUQT8523dB99JsTiS7+3rrLA5Y1HXCBqpKXNVTwnr8t1R/8ZU2vvqR
Z+peNGMd4t04Hy7V5/JHWrWijeI8efdF4V3TPd/0p4nWGQaF9zjjyUS18XFXDG0v
k61ScTZcBhyz3gzjhfJBR0Hb+HMrC5WPvqVenACcaeGYndDv09ezPczfHqYtvM1e
ZcK0WC6VlZpbrEKbsHqrmuesr8OnQNBXIUfbZH0cDnN57eRETgIvGfThY9GayHCM
+ocYB8V5H0wtmelGnLynxAkbfVNGz/ElSiwBM/7H0S9uJ+FwfIUyDxiK3SisEHug
TfYSm72qRHWnjQGFSuXiewD1yoTM9UZaTcSpbY8HPZVok3yZwUPDyomjYA9TGqWs
L97tdA2bItld/NTsREVlYBBzOhDIN2UwgeWutE7EnDvHH3YaJz3xE107LFTh1teZ
I/5gNSMnL+DZobRZV5zQhOUYbT3ai8MeY0o1g06eUAe7FTy1iBJdSKV1tZHHd/FX
3F8eIdYFHJgqn+X7H8pvseN2RuFYO4arQcjCnJb9+3und2HBVVqMZQ5mEyjthsW8
AmmzsoSClJe9Gjgp5oxmb+8l7nGSD1LjbXOXIWLZ0pok+MioFtlzNw/JlJW0kcM/
E48MH9PzeEd8IZ4my+HZpfJsrLBSLPDL1zLbKqnyKFYuieT/uEfP+a43rrTeSagQ
LeUZ9KGeTOAZpVrgOKSbj9reHh05nqvPGvDoSfBN+6ulrq/R3gF9MRmieRve/P5y
5+UgyfRn2qVg5ltYvD9ZBMOJtdeNu7T+qnQzDsjAgWCRLIbbHEsWDg+XkNWKf1dv
tkfwS6KIudX7nu+YUCsu1DbtppNxrHdsq8vL8UTkpYsHn1/U9CiX8RyJg64hN5t8
19Lds3DSIgTVI+4KwKZT0SicMPKnmZ854fLZAdX4dSjvqr9rXoUmPP5t8Od959tq
TX96lwcquZ+wywsJEkvS7bmmlkTXgGe6MRaZ220jdCd/pueMwRN2QWxEaTpFspg/
ViNc0kT8kH5D3Sju6RLd0bsR41rcW5ahciwhj5tX3i7MGgB3BSRKghlR3LqzeEqv
edNbMC0438NUK6SvG2LB8xvOjWpKvPeUiXHqfmtEROR4g0jJvd0Hp8Skm2Abo5qu
cIdKPaKZWb9HblAP66oiUP6N+YdayrgR2TMWma9i8FmgEmBpnWQCNc3Sdv21XuPF
qX5e6uLcvQvHtVs5ZLNSY4bKdxDyVfaT0s4NwS+HLqu5QWQEhz+tkmGj9f0mdgD7
F8QcWAWycQw3FWY4gWWRaQfajB77Nwx7sl/p3U+lVGLGJlBxSavnXqmi7RAxTstT
YW4Bq4qcSU8JcHhZVMuNe1bJR+0EySnhOuDRhm4e8YCy1dBfi7Q6diNJB79LOiAo
7avrpS8l8Xytvv0KR9T6MBLyT/m0LG6KyxLw/kfPBpct+7gNko2TpHFuUghfxE66
5W6ftyUYfCcPxkjX7id74PoV73cK0Y1dDHhY1rqw+puyre8m78VUsSKomGc1bmGH
YYB/Oq+WzAFabpcDpA9mlsDmTqKfVqmK6e6qlZxG3i3XzkftJP05jtsuAlWxSCTG
I/4Gcp4HEGF3Ec6ilgWYcDoonwcNlSTk+faYaSHi5P05TS8qwHctsAngQURz6Ovh
sbq+6CQKgyqP/H0w4z134lRts19rqoX463bmntTUu3bt57GizjD55M448mmsAghm
LJfrOvKxOA4hWwiUnhkXu1OIxzf+5KwD9jk4bv9uzsH6ZCQHXslbreKNyAYNJ0hm
ZfRDx84HykzWiQcDj2TVBeZ5kUAbYLxuiCB1IRHSTYBha4Cen53Pq2VCWOXeDDUM
Jpj6L97htRNxV+Md0sOf5AZ+vuLyWUbPWQcrLqUlZeUPqupPTgyTxC6UEd8xc88l
mMawPr/iLh7FYPLJ+wzgzu76D7b5PjbRMh3mZKSDscZ9+xVYdgiXESzq0G7OTukh
Mh8zpFiwD197kXnrD+wFETRXNZ8KtzXkSLxZhqZ89iuQQb85rc08OypSkYjWSmAt
fcL0LQAce6KJNvgsCTpbhTQj7cF2yeCUMr01uV0jSgPWPGIlvB9VKhFMZRRg6a+H
20hE+s/uz/hPx9SO4Wk3YRNraGgW7xfX0hcyNOIIozqGN/etUFLtxDfz+oo8g8AT
hgBl4xTnQzjOMY7Ui7oecCVyYiEBTC40dOtBf+rbuSNbTKAJpZGSOiE8XUCO7YQ5
dpXohSJKi7FOAmKObl8T54mC0DiVCFWKaHGYr7ayp4pqewW0HkYwKdioFQrmMiFV
SCu4gh0vUbUXrrp8GjuggOVV73hnaSeVgtADVRlXcvWQDEsN/msb07wsn/TI4OnK
vI9EhXBzbD/cpfY0oHyGHGuk13Xo36gpJFrUSsqeAGhHh30o/Em/W06JT5C9KM0p
6X3UQq4M4dKYD+dxMkbK+yn7zREHz+K/lfxk0AZuYOPGh5qIQmMHnG/EG9LHicC1
gyb6WmY8u84Uh2ye7FrqV+/hC1HvgKw7TfbVOvYaqce5h4TxZmiR/GeqijghtADm
DV5cgs0YX7ikRgKpQyDGXc+ezVbtE6HIvE13+TD94B8aZtLWY0PjuTTjiW78LK80
hvgoxwfi+G8ImM749Kxs7DmyTkQInHrChCnrAd33HtxTbY1axO64qhSySn2B6mM3
THqFbQWwmy/fgHetzUngRPM713i73Fi1d41uL9Iz7kjf+lnSaSe58asutWHt9y9G
9sM+mnPT8pizU8LeumdCOeyODcK1l2kOSExO/k3ZBFe92oTHpnAuTsWsad/AQhXo
KkEUEChQEPQ5Js0mo7M14yujJgDhMnnF7HnWxHHV598A5yI/7wPEsurNa49udbjE
0LfK4GTcusWUXdG+dcI9XtavXnlMZbbpQaMBHUpvPTI=
`protect END_PROTECTED
