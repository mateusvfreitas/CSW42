`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FPDNrSSixopWz4GyE4uN/Yzxuovth+jsa6++LQy7r6dLvk7HM6hB2f7fPMQCT5ie
h/lYYz145501avfbfMlWzvo460UkaU90pPzbuawSQ7YUuJel5YB6X0oxeX//FL8g
VRFa4UQekEKAskreuT4KrOOZ08IheN5LhN/iYMYFwyERfFD/PSMZSYNmKIduzQj8
bWLl8Ln+YUtKH3eg0SaADntiifPSlWuB0e+PVfyptey+D96hCo3s87+YJP1hQJAn
G/krdvH7amL4duqnjXjD1imI8ue5nyZfwno2ZvKkjBK/aP012tb+HzV/QI4LDCwJ
1HnvZvUuFYEqLBEu4VrQCwFU8KWaJAJ/s2kOcWpAepeKjc3EUzBq6yUHH0te4A5A
9CTzXijEDBve89M8Q4OP60Mq4m2DqCPOZbPBCRQ+5ufhiFaII3GTcFcD82Ifscab
UonzLyPK7Q+CwjkXnfP4cj4WpOKUErdhkMqj+xlwHwYB9ZdhzpKFcQPn5ORaFfJo
q47jCGNyEFTG+cXJA9x3ePHGKu/5su7Ltc4hrZj88J38HJQz0TKZoAm/gqjrSN3x
SxVcKv3qkjoD1f3FRsKbLd5LC2R2ouaF3qHRVfIEDowL98y7VSG5k81Sl0QZvw1c
0Ptu1VQ1V/BEz0aW1nPg8bQR7qEmJVvyKzLgaRbpzh2TVaQKpLBqHpKCf+mvbRjv
ZuX+tvnEf6X152yeenSy3DS345X3kJDColeQBogZyRrKG2p6FVO9sN6rpyITiY4i
GvCCm4OT9Tu5bDHgyg/iEXJ1cQFCGTFVF+G4ql+aOeUjDHDfB8Zu6rX2P4/jV2tu
Q0JUHgxQ2z/896cYJNhiR4Nb+c/Z0AGdE2c1p6DufHx7V93KUbdhUozkljO09AKw
wk8E3fotp8Rla+fCsodVgygybcB4BkV5fXhXaqAxRTlHotcBepvk2PqWCdDI7R/i
CKDLp/gO0dOzlMQbHfR6bRxDBdzngZc0hAa7ZGhuGDFXq13X2JfdpbDJtoQYa2Y9
+mP8ePdYM1UimeMffr49ymZrEH0eaAU1BQ4ShowFA/CFqimPQ6vOHLFn6xvoM/HH
m6kBBFAR5/dVGSrmkJpoGE6kkP+EkrpqSwovE2PHiCij1vVjQDhH9/NI+Ub/PUIJ
r0XHMvk/zZzLnpW/zjf8fIqmHWauYNmk1ayEG1CgDihjQiWHzgrmSYef62xctH0n
yLrYWKcSbI2FVIBU0e/4TTs2MWXIaodr3gofw6I+g7d3S6etWARAtsitf5PF0d3n
CN6HFT/txkgks0Gon1uVNeU1Pf1xnLmqN7ZiEuJZcGFpaUMcDUdOGi+N19hHeGEe
4WsCO7UBfevMj66uGSJ9/1xkzGbtowHfkXzwELlGo9Iy65pwNwKExkwB94sOYjRH
9cArjqZ6Ie8WTYSA3nJaiYsEh1oCracB2FMZO0tBNKixAgVMC7dbDrgwqQLzWkMD
f3FmRtW5SMjzSyQ6+mMzLppbmL45tjbpBWbE+DFauCQFiizCSLjLOTYZWGHBtaYh
Wwm5IuWyjBTjSuYCtgm/b49crRkt0nKjrXi7BihbYxt2dk/IhomN1ePJ4YpeM2aV
Sfwm2evFuiyvrvwtu1OIFy5w7lK2Z/iEA60Em86wrndGR5378O3/3b00eBZIN7o0
LcrppWzkbcC87nZNcf21vWJyX9ETCSuMCWTlxD4gkPV2gpXCdueTXPjbBoUg6NN4
OzQzV/M1gZMoO+a55xhzRZpPBWFIhXiyyzvltYJ3UcoGso6XxGAi7sCz6S2ieoS+
4XYHhuoeFJFvEHZgIFPsP5ijWzd+oTT0jwxEL9SgG5HYqprXw1TiXte3yhA0FzZW
RMDl3ffwrEh1qWNNSSv/2jATvD2jBm6jd2X9dbWxzyIULcV8wDcvmEkoYBi/6B7/
yywK/aQuJMBB6i8sZInqq1UJVWnwFT28jBEbjz4zryxNR83ChqbT/KySgP2v+HZN
xVti7ZYP1WiBcBvm7+tNhCui2rEmEIH3gILDBcxYFk2hDy36F8uz+GSz5iEy5XuZ
rEp/NS2D0ZClmRfT9QwaZDdNzTZrkyUZRXJYZvvALEryYSTrcxvFVF5XRVu9aYIm
tyxnVtdAGWcrHtmLo8N6OahLu4BQRuGxkxpsXiRK6vS6jEVSleYAzTWh4W5hXwvG
gTUt9ibP+lSR0zYyQCyPXa4ABWuKs5D7BSLOZClM/HuGM6iuGFnpwfJeHPQToXwq
0ElrjLdYpP+xZnEW4/g89g==
`protect END_PROTECTED
