`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qJZyiOoVUz4suI1FltEq4KI67j5mBWVyMOkalBFrS1V9BEM4PR+yS/hDDrnr+rjt
Kao0hx9027kAf72q1pYtkGj7S2dV3VwWK+R+o9480O6+gJszYpcuA8cSbA9JXLKm
ie4qxN73mWagIwd2cumDN9ZY+ix9Gsg4TkDP/yPMLvgdv1s960ZIXWauTxNaDZuM
ncK5m4iUcthwnsDKT4SCTniJM+QqhUGX2qGgJQO+4fwTAYP+8x7RuZ0hq9xMQDyg
G/wJ6rL9G6WQ8rUoRCbmVnwgJK+ZPghUhpPa4HhjygzbK3bv2VyHBnTWiiLEdbew
q375LXwkg4n8o3erKG1iY0tjSVvv/Z8ptLRt4uBFn05HKyf6d7oT3ZkxtHCxBQC1
+G5rShHZIBfv6xCfIngEd4CJsiB6jY+qHj2xmbnpF2QtRPVyxoC/iV73We+b5QPc
RgqI4Os5gxvrbjNNV/7251FT4BAS88lrdi/ob49sipm4zi6OG+qrWDu8FHaVE/l6
sgbzTk30qTlVdabfM/C7J5tG1skCC/S8HtF7ztPoGhnoylcw3CrpY4CD5up28iPm
ylSWAORfDAz7IBp9kGYK7DNH0SbG2W51Sm0EmV0a8yDPxQ9hFqg3FvKYeQJwkiS/
35qhhI07KYm9caKPMSxNM7a6XXJi/qhknK1Wc5j/Dzsz5122dHhz80t5VMmyTk8Z
HIhI8rYB1hx7nHqhOZHvqsLqXdDa+Agx/MEvKJdTkrttZeyfZtYeuVgc6RYgjkc0
xnPKPVYwSZujmtFEglKSYSFWB9bQD1I9NAr30u0VBbmVH/e2mHhTbNRUdxMhvaOP
mKrL3UTB4OJOxDjXW4RE96+PCWsqwwINKovIIQ3whpyjaMCZpBoZ3X5/zrLs5M5a
GagdYpGrTsgxlXKQ9WngIW0EIQBx/RCwL5QoydlIas9gRv3+qo2XlkanJeeZ0lxY
8gBuw227G/RbGmfXt+uoUt0kf1j2XjMRCkOASpeXPtVOtrEwdD6gLQtSD+xPWoVW
QLfqtfOQcVrKMWENUbbUvP79imjXWOOtwv0m9WUGeHXf+b5KoYOKRTdbWCxBAhEA
Cw37uDqAhAwn3bNgC6wR1TtR6li/0ZLdJNhk/h5PELJ/NwPMrhKHfbO29oWt2hSe
OdclA7tm6Re5Xs9yVBZeo5mD6jOuIIOIXJ7+AuKm4/b3BxHoiL0Ikvb3MKsI++ft
1quuSlXAZQ97y+x4tpZUS6lNvb/frrFpN3YR0lqJKrmZFoetfkCxc4zsMJ0QljDy
YBA94DFB9I/mLdZ0sEhegylXjlbVcR0vtYtXiYQ5Bv7PCKl9FXnkXhbOcAFYz2Zt
3KzlX7CAzY/vT5244o0Fhgab7n3bMYMri1PMlFEiCi30scEmOj74sxnPA0mM1Kn8
PehQIUOUadILOu9STwunOCJP8AHUBSpkZH0I2CkJ4cve1s07RNl9ULNANlLMotWm
haOc1dQMIlzBDOFcUwEdMy4UJeZ/fpJvPAfGlrvSNuN4rJCjEInYkXUdbcGb96Gx
IFtKVBUOJwUthX6oxA5nLK1YpYGA5a8qavS1ZzRcVlrifkEbYpKRSdP4aJ+40TJH
Df8+RDBVku79e+U3nerIvt5XLaJmtuaiULkhH08hjCfXkawogcx6sYl1JAWBqyHI
IXYTfas+G9chrJ0Kx+OpE/Bm7KUzWXY/Lfhi3FQrgI0jEWPb6iGDwylUeCZHEGtl
xN8iU0VdOvCoEZ11zzF2gSpJvnbjbaA0intYzIzGE5RtrxRz+rJVI3+fr+Bfmsr6
cR4I7iw6HUIo3UhEzYidJhOtVJhjtN84j28ts3yh5WyhVEPcAnr/Z0p9DpyBKY+Z
piV/wDJznaji68YODVjtmH6ukz0co0zm5IrAViFBJqcqU+D81SfSiqemfOhksgTZ
SkPVZBUxjV1DdkzaLui28jd8PFjuifxhvPS5fGakiY6nyrH7LFS7NdkJd2etg5QL
x6JSgmQq9AdEUZep9M4dKTbkduI30E2yR6EGei//YtTGHWkAzkyVgyl9G2MMJKMz
P15D5jyzjHC122aF7xFF/f0GLL9/07NfXz8XP4ZcUlj0VkBmURdTQixz/xh+QdNn
6f5LYYn25l6zNyp1U9C2SWapo2H46s9HcUgZ1zZEixe/GaLFa6bU713QmmETuOUK
6Wr1qGhJeRRGaY11ogd8Jna5P4qUI19ehRMycrNheLPFAOCko41uQGu6PUO8d1FV
QiCU428oPboEU3jKfHZy2bddCGih6kTuioI0RZ/lhS3jCkqf1u+QY0pRYIqktQq9
pCnQscjwctle8SIGVEEaZFBkTf8GqEfzN1ynJdKOqXT1MtMxsqeJ9KzULYuVlwFT
FtXJiaDYKqG6e8aENbq4miOQWypCA9rwLYfI3aRD93/4BmMcOVsS0KNfI1R5/BII
coBOKc0P8AMWJOij1ARYV2rXYidzjDZ5o/M3D1VWp7zQw8kCNASQQv/SrSzTddbK
ki5WtZVb4v2EUwqeQk0kOUF+e+F9ExifokR9jMJyMzI8VIbF9XgNQFfWCNj73VcP
2xWGiOBN3KQgNpornvaAVYuUgCd3H46PV+ktl5rAWq1XCEMz9Ady80jngPzgUhiN
nSpDPye9Y1I2UEmcayypSI7vAlKz69XZfVm8Cw0/918UGGf0Bdg/DLq6/v24esqY
09zwyR3/dm0K8+TqPJsAU9rOaCmjePBxNP/a3JrZhg9PNu0Yc963lzxbn9CemGKt
dKgL8AJOkAH8vaaOmew2f+R3dYoNCutreJHLxFoKMI4OSh7mP8P/Mp3OgM6YiYmU
iu1OVmxzVzSRs8e7px+hho4UdKciQ1c/usySxObfvcjPs3gjC71yzF8XPuKAVdwX
p55UWVFfz5neqcAjcA8xgsjcgVpkPYAIMWiaqGFMthxLRv5tL+e4KRA6I2jo2yMJ
u7mVGNwh15jcvAsU9cDEPw4UwQKKxvRLkzRSPnKMcr9CytXjHSFJJzZznaYOx5lE
EjUByNwtbc4lgLDujgTbvf2ChuL7VpjZrPRu337U+LU+aD55J1bmaEOwxJr6tYCz
W03CC+KzkxzE+nuFGl2Cn9pjoGY9IJEQAhm+nz8ScWRR6N4DzvyIJa+yO2sgA39l
9AbToD4w5bMqnUyFlxhnYe4+4f/M8i4RmXzuExmww9YawXA18YwYYc4rRVQR47C1
r+g6S4JE4IxrFAwsrQD5+mZAvNaSStQsTiPf/KQExLmhMZoEP8eZeED0udK5areb
r4pIKg0NNefnzYAVFZnQ3Fg4OJRyWLoZVS3hmbVDhCZQeyE7AA2OSB5WUJg6AuR8
9H/An/ureLTxzUi4C2YMZ+Qzxow61KWYIQnWv0czOrf2Qxm1xOcViu2OD7mQA6pA
u7T2mnxkGTj0pgNX9dSke+b2Wb12jZdwVpXEBRyWGSCsGM5RProVxg/tpI253nlO
onc3Ksl8g6IWUSylSxylEDJHxmjvX5zbgb0q+sAggeCgBG5aCwKuRFHvRXVa6Syx
I9vioqZQ21bpIfZh0EDUborR0e4ztsjcYUJ3ZlMLUXnDEqfcdJ8NfQMq+wFRIBll
aTULKN/A2bkx2D+AoGTe5rDcpUS3eXpbITzlkN0eQ3lwcAtpRx1mmDNSyjpxK5qJ
KTMn5a/qJVG+Hx3HoeLdc45W4V1UhVW+YobSxIsI0R+kZ/o81YmeRDvAZ3lPpWFT
/B15rizRx9FeUmywtsHVmNPUVBkL94pu4RrbI26nr+VmOtkBHQn9l66j5semSB72
QTvrEFTraP9DdUbKSx4b381AhPngGT3LvVvEav0mDIST0vSpfdCPEsxsMu1zXDKE
CHO5H60yKk5obGBizdMjuL0uN7LWouR0SQ7uYNYJhd38RJ82rXbFWks2guh5VVz4
NkX0I0itfMfJPeH19F5RYiXrcU8GIBczOdKtDgtaLdZRA+7PAF9TJMiO7PCo5qXv
HvnDRAvUM/OwXInlWGa0wd4BKaS54dxDQrbM0GBhM9e4qo70f9Gh9IHGLsJMrbFN
64jj1Z+Kk6MUsy/2hb6YSR1ixSZ6wugS8took0GnjJYbbfSW8J5eP3X5M0q9o6Cc
FY9Q8pqjiHT7tzp8Ry8uyWJ87ajOeXmya4GBSCGmYS4MvrlW1EJ3Dxdegd4p1fuO
q8q5vlHBuOIFs9WlUfLOfNl3fl/fMjtHlwl/7RVKK2/yRH/Y1Dw+FR1Ov4IbSlJF
9UHviMvyjASi4PJygigtAkAvZPEn2d0xUIH/AlNT6+1moGB05Qk4NwB92ro0ne3/
IABXcCoVJjO9kMGO6D+IdEUoMwqOVTP3hsw55NUQ5jvdXxvQLfuQQrMBdqGREUjP
ogpOg+TRk7JTRYfnsqjsOg5tvhESICA0HmPx2t4UyBiTt/Y0CzR/YAwWV5BzxmpM
UcTGeP2BuAyEbq8XcvqHIA40kdxjZvu9Boxi0b6dbDNOoPiHr+Jscg8XzphPQf3X
qT5BhyQqVQB894bbI3hiybhJvR9t7JpcKN63MlKGy7bTHgZbeSuiut30uk94w/34
iB+5naWQwORugaO/wDEiQCeLQ+a9UjRWQinKqeeCpkbumoCvaxwQkw3WwElswwwX
F8GZ7UBqVooBwTku5MpxjGGMaRZYVForZ5ekRVENFY98wV+uHqBU0uJwltdX56Xj
bZEViQOafglnH2VdPuOMJj2qQdqq1MJIzgrQuzGgkIVTEXNio9mowf58zlfKvNnz
aMUBNDgPRpClhaz+0GIP1r0BbvQb1IQYQ1bIxrruA2zzqWD2Kr9SVHDyWS2JH/yF
QLOac37iC1fA2v2Wu4vqjEPKaVcDibqe9T5ER/AJT49APFwsoL3hfEZh3vdSAwPe
P5HwkN5MDStUqxFbTN+ig7SQTeuMoXc1oYA+HOyrgDhjXRN6ZBZdrGK2IAcxrLJH
htYn0P4OX7ineY4E0cgTZ+d915FvDIwRI6wG4kTLvT6ddGQ/CXuIO4+gQHU8iEsQ
PhdjU9Sx92s7k8U+gt23QjC1k96s8Gz1Y3QJ/YHmbB2qIR0ZTjwJ9e4fR1vn1Rt0
V0kD0bku1X6+sCe+DYb9yCmwMuTtiAG9slqUB769ZHX8H211QFJUBiVc8KZo6hqo
YcIjgFiEI/lxAODA7kr8rJLlIxA2oAgj/KVrI6QfvZiH0XFcvpfZUBCMlnUd9f5T
gKgyOLdTzBowrezikioVbc1T+Kfs2g+kYVhN39prjTXox5rPCzpwaf/bV93mPvhB
/zvhJigyfcI7yIi6YR/wtsTXwiT4ebZXUpiwEMlgkSTxQJMwFORQd4/U2CQNnX9s
2eT9HrWoIjmHd/IAtFaINWBApPdCJBI1j4R3AWsKpFittV/I5siiMNNh/CMVU3BG
phIl0wTFKTmPUaSK5QUSw93MpmaL0AhLqyrem4a0bm1PdZaYPblj967+1OVQAnVr
OnLk3rULHSOPRbGwIGckVkFpzlRgkW2qAGDdnU/2HYKjLdM6cFsB7dkUL8eRK76R
N8w9iVogDmYJAGKhIuMs0BjxVKoZrLwZY+dd8qBH54Lk6jp1aeSBO46S56Xat1te
OWY3bXB7G6R11JTa7bYetZ/r42uK5jxxwPd8maLSBkSE+Dt2hypMRTQF8+aryjV2
CPdqbpi4x+IEFJPkoyVreEzv78E0ATtlg6G4ujh/jaTwKK1WcR1d90QIj2+y+o3S
T/SIwzf70SM92m0TIj8wPEYgJ8NFX9MCNpttsU1cehnkwjv4DS19KWr/szYwkPWf
n0nObvwvk+E93fOzXzlkH4VZAlvOHexld+6WOVqTZKluhnUUo6vb70nrsVe61JnL
zqd6iEphrvoaRMCA0SbXFwx/pi+TpVWD6dfr85tpk/w9M9Iyf6sXDsafEmFFDKZk
883KJqvIqx2gJ37as8DLVlJfIjiSHlwOlFjJedZe4LgcdCldbxKSq3pcYfocI9Ke
TU7XCL+bQQimupETCYi3veGFWZl9wsQUgnnq6CRldE1Vhb9j2wvnOO9rK/1ogk+4
k9SXv/lViUWaKV5IKsqC0GKaGK8IFTGiFsoX54JoPF4wp5BBJO+b1ZOUBBUgxQoT
Mf1e0T9w56PwNn9dZG+bxh92asaiSc88IBAWpfQhDaYWvhGT6M9npiEwrh33TPPN
vFTP8lvM80UvtxvYqjDPpupl2cnI2o17mRDRvGApVckA+hMg9rodScrrKCryouyF
E3YdD2qkzvOXtbdanxlluYUf/cPhAt8sVAog9qf9kot/fHMFP+CuaJgtdV11YPyG
Ii7JkKy0Psk5TkS/T0PnKeoxo6PmifU5RGng84uRzHExegGgA17l2qOi1UaJ4naZ
kOxUmD1FykFVj1VvnARiKQLKu4kO0behPGSCq2a73RQzcTMzBz4LVoeH86KZSCAT
YtPkxC+Pk43o7Rk5sRvTP2liG0N5SmgsquLMsx+Cj2F/0UHSlhdKwtatzTEX15Gt
3uJoruQlKNHm1z43p+i4Se1MuI7Ig6qsotJoBQ2Yedt3mi6fiZJA7+Nv7+3W9xaF
S0/G+g78bjwEREpLp00Rwu/V/5dgTxCxrRdQiVDkn3Zd/jXuKnUDzH1CDt6gopvR
IeiLyo8TEude51TkaBxVD3uK76fIACQ/R+jejI6YdJmXT6bG51nRax/ULcjxVPwd
rmAiyzs4a804HCb1UDa6/Spq6D+F1ifQc84t/nv/bZsQOLmxhYnijbKaVm9GiPuC
L/WkQGQExfc37RGHrevALRccybc9FqaxpQbfTn/45x/DtInfOBdXUfqPaJf6Gd65
itF/39xjYbQzDW1d6p28mPgqAqokwhF1LOsRpDN4BhFae7eMckYcEzW218p3cgLw
PQ9hwBhj7CAY1gqZGRctPdCcGwE0vYH345o0aEcCiSJRCcyhIJl7JAomPD56ShDc
XDwzuvOpgL6DVMZB/34kMWm3Ym7CVhz7Z8Snj3yZwJI1IXn8NjK7ChDQ2lpybpqQ
LV8SBU5GBIy1xl8e15+nrP+bRidhXzcpVz9f0qxkEi/aydtjjDx9DBaRf+PGnKcN
eldxTlyXN//tloSQMou2tV9/Jd4oHycdEf/HRIh85Uu9tZaGOx0CF/9EhIWCRfTm
KQp6HYpXKqXRRVTVMMxMbWiCogEiKvNFii4QrG593iNbl957bpYTEDn/tUbwsF2P
XX4x6jMjGZdMheFGNd/DbK0R/C3Il/2pnAcSpihI0KzjgKaTECH/FoE943v6HvX1
ZN7HeOy1u9/jLv3u80OnS2uJ3KZ2k9iJ8WykdXM0GkUVVa8uQgPVraqlJkj0FSq9
HSYgIP3UE9c7PQpDMf/PyRkCOQMIFlR3IOmUuGYzBp5oj4hQGXMh95tL1PCwpeNN
8YV3Rm5wZxebThn1rvg+eh/v4M8ZOi6BnYgyaCxlv6wszGc08dJe/O3fXLEtlg+o
wKpmlrouTH7M1KquWpucOsdMOZttrn24VY3d2Ijv6x7+Te2xlwCQ0+AVkQxcIMQc
DJQQe8zJOFrxCBCzvpJZYWzbT44oBuHNUdAeJIcZo3q1cB/ziH2gRzYmnTmCqi7d
pR1TB+4+5yc8KJtH5rYBD4Kw5Aqeldqg9F9vD3KfbPXy6oKCGhrGDfq7tZ8ifKY2
1TEi+WKcBIEaMLegq/fsViAgI7yAQITeqTCKvQqG+yMHFHGQHfGTh5YwC+VU7meT
2xKMGZIz3A3HWdxFhuEEmvcVTANuxEnigJAbJmPdM7s+Eg1fIEqhE5GdMU7k5VSN
KsdsFE3C+6s+bXgykeqBuY1UyNvC71bL7/H/lsVZdn7Y5sA3+K9K7ouEXpZagXsQ
fCGf2xBNO7aNZ4jpJrb+uueo66ap36Q8y/xOAqtSt8rWjuYoFNeIOIphYfG85ky3
izqChoIthM2bsvfXxEvB0OyD4Otxj86lJgG8KoJJ7ifdMCYKKWCf9j/ccw7cOApd
JeXEcwVhCgy5nFvWR1EMR/5sLjETdz/TD0dHodQupyHY5VVe2xTB61U6rGG4Pl21
qhkql79QQrKhFxM8AFnAHBBkWSnWhjJJAo/voWqAMagd2uIqeA2K8VhAQvP30uAM
KTajF1vabUAbd3X9eoYmLftNUeXsjBS29x3xBzvjw9YEhYo3smX9np0KDOUxWlYm
XUYFZSd5Yl8tMFSD6Sjc8tiQGq7DpxAI/MbemuPrP3FtKbelM1+OwSP1CPUbTKxm
wgXkOF727WqDM7rug39V+Ti7f/bHPq7zHImgTHsdVr8QURaXXP59pBlFW02H3nI2
JNhpgF4vbX35Ne5NH+74GyHKqmAQkxFk6hkxSmTQQCG3JqbBI/hB5dl6x5CYz+pZ
IcmwpIZRyZ1RPTKnvxLl1lXGCSoftI6T/XOh8dPAQi7/5KoHMr5PiqY9ZgpkqveH
YRfjjR7dnEWhnpf73JE2WABZdeYdhayHaCL/l37uTM6T1Dqz2X7dyhO1uqwO5MXa
dPT4CXy1Ug6HXGOQ0GB4DxJ+NOH5QMkSCvKk+n0zO7k+6lHw+zMPJ7iMMDz3K4ni
SxM1DW4cCazKh60NCRqKb2im5EfslInhBofTmsDBbJkaAW8++Upta2LdtrGVkxmf
NOhItV1TfrT1TNCM5b1dCEKXgjAzVK7g4fX/OmylgHQmd1WcjXHLqJbnofNN+xnb
MrrH0eq1Vko4YdwSuBI5XKpplGBDEgUjejzY5J2V6INVzViaewDqys0I4lpWFLFV
//BNKEsk9IWv4xOZDyaDqik61VM43refiVZ/V08RNe6aQdLxcv9RuJV50TzWugbA
jbseskky7RdCB+b6MFbx/0RgSuNRuKL9DgcLV0N/sjPm4K5dMnsi2mQffFsqv1ND
22nitMXL7O4AWORwZgjks+ZreptQ1LUJO/LOqw+ntbPscwU1waIE1s07XtOdb+0u
yChFq8YsLBB9/A+iny2i+gtc01bCh/PG8dPMrmaVSq4=
`protect END_PROTECTED
