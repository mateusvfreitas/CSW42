`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Y42LYcAj75JONtKdS2NG1vngP3ymoxAvONMBMlW2OSCiYVYmPzA8ijvKVmWS1BTF
nVtjJKSi8A5Q/dWVc73mQdmrZD3d3roUmumiSfK4KQOkbQQkTiy+YjK4Nl3aExon
afP1aGksspY8nJEkp0CtFecOXLrUlsT1HxEe9B9HGI9VxHb3lgXkX6Yzm9RKK+Aa
9xGTCykFD2XV/oZEWRs1zAzPUlphmutdPyVvwmMUIPnx/nFu+a+AzCdoGqCu7iE5
MDoWt4Nf+zaOlEZqSKCbt//FZtCuogcO2Hzl/feZ46KCUBeRMe4Z2Rntf7i/lJvv
cCoG3xak3hiTEMASRQPV05lfdlHfrxjCLHYx2MDu/lldLiM7NqaUDPEBaUdaz0pk
wbWrgSQqaigU/a77QnW1FqkWU12rxogMIPU96lrtSDbnYu1Q8Ea0GvnfNubKNoD6
BulIDFDipUp0Q4wOKgcGApxuSSVF92AFS7sJnm36yIgAm0TUnz2mSh3q8wisTALF
yTgX8ahBe3rGHs9ot5xEFBvPMOC41cWcavRoXGxiJe+SCEQXHMSxcCa8tuPG6h1Q
jt2l4jWUCwaJfBHTh+n2SWgDOFWhwvz261n0/5SAsGw57SMoQ4OXPZOKIWax9jzE
M6FOFvSIfmvyJFyXboSXTuKQDtJ8du5UMA/fZORd1hApftI17gsHS7Khf2ddBvRt
k9SidAGBU8Kfgn/ZFuwiXk8mna3sbQZRlhyvOfpQAwX2wRGEzeIDDMAkDjI6YG3P
8eveU7zKjiub3eHfq/22uA3Y0fnXXUU+w866ai4Cl2l9Wao/dvJhR63UB6xVvDTE
epgG+6tMV+L7SQEwAAMvw7WJFPL2dgD8znni2oKNmH1aoIbHNj9rgD3CpHq8mz/C
gOTgMCHuHSyI0IOOut0v1l+K6Cj7ZUGx6vOBfahh50PABU47M7rqDafyEF7g92+D
e2c0uhTD3rwLg9YIJ8ixFO2No0JkoxqDFwnn67OniUGEdDRIU2YmfwbrXYfVkOxM
zvWBTqDwL7l1E+w7/2YKW16jqInBuWRmvl0VWZ0PB6MBv9f0OeKoAyjU5F8+fta7
GNADuEeImrJDzUo40EdNwKGm6srFucbX81VIK8Op0oDe9oO4J7tWcJ8KcM997agj
5hDxJIFfSmO0MDeDzz4jegfJv0ouFyiIfVHdr/ZT1GD8g45LKwEgy4qveBooKzdz
uzwgi0Nx19pyHzSL6OCIAytjEsK3PZfrCkpEedy/AvviaJhbXefaPHnKQG/hWplB
hyBAgWP7nGfrv2ARtuiEgqrJBhxO4D4md1geHzn07pMje2Z+2a7MwFJD4IbwPA10
FkpiTXwtLyAgGWw9MyG+Xb5XM0o65jLrwLamsTCfW3vrT4Bs5BNbw3UbbZ2bgW/7
y2zv4uDDv8n5GTnVL4toIwsQmzgnvV9jNDQcVSaW3VvncyNosAEkJx7Y+jZ5WdY6
QmjTXvXhOJzusnXzrwzIagQWVRMSunSnV/vhQ8YCldUPWamNrQWHyNAmiH6KyWNT
d3WB9Ug/jPWLDU3zTGlGj90pTn4zU3lmGqzp85mwr9p+coewvLsYFJ3LRc38vc6E
h6G8lTcunbzDenPiO2oAoXpJ/F5iPFk0nj1nnyTmSeEGEjcZn0BNRpbm88odX6tD
NiONGOW05GEcicYHCKqQPSTswx6O1l6ej4YPAk3CZv4Pr1aXhW15Fus1mGPtlVga
voMMEALkMd84zOykdElHqcIMmyNwXI8GdoTKnHNrbBJ3taXvpQ5hae9d03Chpsfd
S9xQdjDewWkvSEqguMP+U+Ev0a2Ey0eYskwdtNFkLcpX2z7n/lNeCSUlFsXR83AZ
iCtt6mP5F8duiBltHpjh9LDGI7fkWp4DRRMDnq8bijpR+l69cMQkbIyO6DN6rBH9
efwjLb5HQ3N8euwrLFEkdFT3qHsAddjPNaOzF8c8u/lwMegXRPekfD4bYMNSBElm
8GsBWsDbtlUzZyfijLrUPA==
`protect END_PROTECTED
