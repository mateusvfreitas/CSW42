`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DfwkdywCMXg3bW5Ywt5xqLXY253hakW2r61DH3bq/riUM4oi76Ww/8nMDzutbNaw
w1OOnCEqpdSjkdtaSCFPWKQpwrjdDbkErcTd/bf6314DxY3ZMvdTF/zsptn4teYT
Tt6IPxp9JMElW3HKxBtBsDGy1cQDnauGnnEo/uhTr/ZA2VU2KAuW3ReksulZFaor
TdWaReJUl3LXplqjNzb0QLoho86wKRpeBH0X38oDeD7gukK9dzKFqrxaWToDhQsA
+FFBPBFb7HnLOd6E10jkfSugfKqoFaiMaVEfqTzsg2rIZRSPFF9n/JL6oixR32xe
4TDgj5odywcTgtABzBv/5MYeJ2sX9YkrYFAkZ8jshQLuEYH4RmfcsUluYoAr06Z1
YHlZkbVNQG2RGunR7s5YxIGwUKPDfcdkn/gMuClDWy2y2m1lof3D/x0duTptkoDR
tdkibVpsPZXGIFYtPc8xqupwygc+f8XCz8aviUPEhrABL4PTStYzPM1CQkMv8GBu
g6WoGSnoOIJbDN0CSlH4q3soWpuxI+XYZD1gH+2VmnIYuGRT6vc9PLKHq4Yp1vcm
/j7CH8aUvgDtu/jaJ9FDl1NPSxkOXfDZejvqo3yeH4doXgA3dcoG2WT1HrGxF6Ud
wIsQoWRxdU91DomUEWP+tR7xEzRkZuIAEbS6++CLmX5Cly1uglxt2pEZsLfVhT4t
NTpklkfaiD2moZtQQQ5K3py79rM38SXGoZTa8VjbQoQKhsLJ21SDClhqklUu2dgP
lGiFXwZZIz+kmguVvPyRTTqQEP49kNYoHiBcFcW32IuHVXAS9bV8JjpuT0xSdntP
CDWg4GOYx7LIB4AK6JI6Vab4vXKuyVVOSDa2WcA9OVcxGsrH/GibINnMQUCYdmSC
2pZtAAzYbiDGW1i2FgEHfxDHKqQwzzN5Vlz5xwLsMW+XKL0PpYnL/lbzozPPVrCG
WVhoTLbCPuIiOjBPGes8hMpgiOADr4nNEKHYp7FhzvX9ha2OiNvCuyZJ+bfDhvN3
p6LPMl07PTALWLPCbJmjd7ZbChA7iLG8bJaFbRYLF+jgihEXq4Pzy6Li/7u/XLPH
qK8lZF3lUtBti8q8rX+4k8Wt485NfKe2/02CemX9kmEntWIVMxsc65/JS4+c/b2U
2QrgdUho1xMGC0yWyKBw/4KwNVzt4l0yxETgRrTJuCgrhVpP8sqH8unksAj/sQfe
ZaqCfBzChdLgC6w5owvYIXV7SgPDFZXkrkVzGfAJqRoKDO8B9n9TEnnXpUz7xqbz
E9iZm3gQvOvYe0w/27X7Tuht2wtDmpc7ue3TEdiPcsJ+QdBABo5XSon4dwVhKIdz
Sgxv6iTH6zya6lTQXrSn3kyEBgNgVru0xHaqOP0uffVEsWnr06iySo77CDxJbXs7
F4WFx/gZC4uhvI41GTRIgQr5NOR8FLR8x2qSb6/9GwPhqJ9wgN3DExRpk7mtBZRb
O5ubBlObCG9WuYIzoyzGLTQlKJDq0oaquwQrf0PGvh+8/XH+Xke6YnN1j0k/OA31
c7tclje+yM6/Mn//j0QRyoxNobRzwWsTGW+WOPnAkAtcZmRS5PZ14svKOGgiMKiU
5ifpN3QDDOXn93dGuw8w6VbN71liB37SyziSiIF4cEfG3+NkoTIWAW8ZX2MPjLmk
8Tw4l5aw8uFAKqJI7TGbH5VxFw8L6CkK01gjem5I413o+0JK8i7GHIDQ96g+RdU6
9V0RLyndtGxgNh0LaNx6eHPG2n4EDZi1z3zp8OnrHGpiJfyrs/NygB+Y1La6w0tm
QM964O/snqW1gn3oGPYYNK/B2eKniEVKqvncQYlu8VeEG3fSWzoLNKhiAcTc4Cgz
/2GWyeahmHKp6gTzfdmCc+npyD8Mh53ientF0E+ElUieSpnPwwAFCelULraa8FrD
ZXcoZKNK3ooAF1Wv2MfuvnL7s7VhIRT0UjKSI1IT4AdOnhyo3Brlhu3rl5WBPRxO
W/TDbXdnCkgS4zBqNoMSDQ==
`protect END_PROTECTED
