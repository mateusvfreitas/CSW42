`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
YpEaVxW39a8i4jmwgKjRtddef+fu7piTugibul7S7HWfTtmIpVUxzbBDMe1BbKwH
CHki7IzBtSXXYNJ3HAWz3JstAtDjCMpYPqfymOKKRNJagDkv+SDGF14BOUPylfht
C3HOEW3ILfitkve1A/31k2NTY4/GI1dLwzRDt6JLmD78JMOESddTH4GhXWMF/FLI
SnLT4lLC4BD35ZHDgEti1M5yVaMCCHvBYHWT0S4fJjUfpLKM+z06lm5N+Bnd1ojH
WgnsnizO7b8Z0gMtFnG1ACGBJApI+cKzcUMMG2lZurT8YX+J33LQk10CTHAVqLvr
bH1uwNXhm3FKBC/vWsoAcRTXRmC8BI2i1syhbXA1Wj3N/fgSrh7oYkOfFHlBZ6NA
l3SEoqRzHdpHgzBR0g+6yW/cvhsrom/61wI/54uLn2As7f2s0fdPD8kNkE7kHpW0
IJ1GBkjMbvZCTQZszarfyKcT4Bcdb4tI+0zyL44Ih2Jx5NedtanNyl6lBsTCoKZJ
D5FgkCjBE7+54/f5I1xq4K/bXqbZdt8NiTyteSg24m59utJ1u8D2GOVzxRC9AOze
Hq+mR7Zt5eKT/GyfBIy9p3aXNU7iMp1gZVnqVMs6A9DhUAXN1zMe0BLJSElPLjzB
+kFH7TSuoEjRltJUKA4lFJZYnkdOJvjxZpKnJJCYVw42r/47qBCILwh4aBSQg9Ch
Iyj+yf8goaaEsTr4K0l0HZsmnoYTEFd40vx4dHRcJSI=
`protect END_PROTECTED
