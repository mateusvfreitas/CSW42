`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gWyndwb7XaECNFuuZT7n8ummRP0ZuQyE7iabr6MvFYp1bnZ7a+2J6+Xi1S/09MWf
gkfbfn+3rG3sV1DvVloaaR/91lorsvpM4VvrTsPT7cSBr19tPgYc0kQMB58xRYr+
0cWCEC6Q5fOfd6P7y1HMFiLaHpHU1Eie/Efjq/w+aGEHtpfgMYnKOqJTyz+J4zgz
S/ne2mHHBjxzL5PakhCX6trezlF5ApUCGhKzzBNX9NmlvJEGF1uS+Sc+PjEulYRW
i4TGlUkzNRf7CLQ8mM4hbFMFi3wOzax58Aey/VujtDZVB+980xBLtbVeWhJTJASa
uA8sN5NdqIJaZjbaqqtHt2GPl2PKBc7YgkAaV+wbXfamDYizPn4Nf4s2cUy0/cad
Zgq+/eeM+JKHABwpC2q2BbfL9n83bvrlLPjcOeeDmyaYdUgxIKHYUbDmy235NhWh
mP/7lAw8YHz7yY5mLn5m22+I1AM9Ueku4A6IMnVUjDRC90gJDpZ0IBziqI+yGu76
Er/dKdg6+tQSiaX6vLXIw3OsWaCECvFVCVLvcyEm96vr2yNLAK/kYd1mbPi3OCWT
dfeVq2nZIzry3scYkqLDk77mwRH9Ndo9VNZAxv0PcgZDaUOWHSSbmF9cM4j8qyAL
hSYp0dmZjLdLJkT5bXEDQT3q+RfBF9KB5hSHImdvhWNw9PcvrWG3/kYJoVZjmug0
1IGYMzx8YNYBt/kvetavYWmMhYiLZvqCqlu6PDI3myyxzL37tozJUVEYyD/AZv10
uzEXCC1ewSywwfi1zn3F2hhlVEIkYWVT4nbiZfWyNSCoByfRHGpsfitznhEGCtnF
JCxY2ySmM49mJPRhbWcK/VYigN/npBQlQNNWUYoSr6Yy87NjGiRVoPcY8GELNvBb
fc8HdAg2uLxyTPTbeRN2ITy2i591I13nTBDl+C9KI2mmNGLEco6dedqjKtP6XyfP
3ClK4sYGAE5DEBA1FbauFr/Xftw/auhFVsU/KLEUsZQUJD/KthO4oZEB48pEwkYb
jK0FVDpYc+z2Y7/uogYzVbexfe6M3cDF4PCvUocm1+etpKg55OiCxLYftIy9leFy
06EBGTvzDenvMDtDQCYnqcEvG5SejXlRu4yI49eP4IKfFzvqpNOhxBdJ105qNQh+
hte08G4Mt8E8Cn9BT9u4PpU5nhTRpmn09/kcPaSObTr6I9ZDEGWFxOcyDFeNEOLf
bLMriZmPAws5eEMXv8vFFkJ9ypPfC1ugl4zgbbSzQT89PY2FnYvYONczHRIN4E7l
fI6klU9iixbAH04Y7QJP5S9dkezeQcnhcI6y7/ZIoBZ6Y+LAdponAbuY6OzaMaKQ
dVupExfX1ayQA+Rv0pSnRijBeCSFxAfG1mVOdIzw138L5Syh7GICG/+ZKQtnJVzp
E/1RGCb424mCkMHBIl6UUJLVCapNgQiz2ktjLALC+PuKA2Cbo4y0Ii9zQXtxLk2K
2eYs7coNyFgAw7uIrE2VaCMNaoeGuZELO6zLb0bWbHTX3WpVZ4PemA2+mCXg6ubi
SsHWXcMsMeFezU3DVutGRspx94pGHrgCPofnCX1d5u1b6uQhKoad8B0GfA0TQe+e
lpEd1z4TvfGTag+KoFgrfj/xKloYPuQ6yN8L02WceNp3l50inixs6dddfo5R1spt
JO/3hG2dy7enofS3qSxZ6wMW35WjQEgZpxiPfK+FnuPiMWeSiEUyNcLyJOezYagA
1mDw93yZcLFDhOUgXEq9IRlpsdcqQBvF93hQmReukP2KCtzEGDMZPfo0qumP8bws
k4uAC+IsbKCQF7/RejFtIKhHN/aFD1qOe0N7Cw7HLjWjkwRRQsT034BNUzmgEnlm
HCdq9GpPacj7Upuv62X6jUWFhvSsMtogBTQQewoZPV4g1Y68uTiznGynMRGmPiXx
Sb8anGTRRQlfhbYxd9r5XNXoxcl6EeiyGGZwRF9eBw4NsVSFiLTOXxRjKL4NRfsz
VzaZPkEqfhlk7QFv4HM3s52w+k3oAAtqEBaAkBnsys1IoYv/jRyI3PDkyZaIzSE6
PZcYmaI07NQr7qvRtLO+Xha+pdkiK16pSz+7dnRtbshthTKLCaRLyYt0r9scJKhm
oC6y3mRqjtFDVzAF90GbI9um2dchOZET9BFupHKvTTE2l/PcqYfSJyRRqPgesz4N
l171lZWMP1BKWfxSQCtznr1iqtDF+7dsiYGUu42gNkD/5hMcxSi5ApzBISqgsWy8
cW9NxJJ3A0vHgMBcT3CgJTAem1tVcbsHBWmSxV1sPFnY8E6IBbtquoeH1SSJGHSJ
JVxWtMQb9zlOQNnsqjTa5T9CvywcqiESm8/ty9ozbroGLnvVupF0SHvLZozua6e/
td5MeKtYER7y4K1DJRgzXYcz+a02dUaBHaPrm7CV7mdCmTpV55qM66mtdUSlqEVY
71zBIMr/HFjbzwig/VobFIGxZQO21LllPxTSxhdcGrKum7O/OFqLxb0MRx3vb7Cj
RHX7dnFLCRgN9P5V9QshXJDlKgVPW4guMZoeWf/jLU6YApqxSK3KRhehJpOXJOqg
ibxjzRUYlf80QPsFsV9snjm3uvNjA/mwlyEp0xrue+zlH6hwqxQvPnYMUWp38pJ+
azxRAbuf+LZNVE6qy7btxikGisQm4hhkWwYjSzp3O331b+/9vQot9xcSEc8eF7RV
bp2GkCnkrSKshmyT/YRTXjAX6Ane0v/21+Mb4+g/DuJaqhr6gcH5rYgH9WODRLs3
TlZGTDk0CG8zw7Rwdnr8/UhDMRsakiCdynVgHOkgSL+/xrw4a/q8BH+tSq6HYq5U
b5+GuZoUSYumF0KwlBpgoy+tlgvPmTrjoFTddTQU3VqI7+I25jUzKo2+8LNY2EC+
M/86mkI8ETiGCRB5sPbrTo6CsFYSvCZno2rcAwDJJ3TNRucj34cMxCHdplCGSS82
X8CusHQyBACI4CVlDcUi9iL9O4ZSKDFz4/fK5YXhpurskF7VOV9GJXPHO7V+928m
vslDM3WGTeh32iO8ySRUwn2LV+qesaBOCfDRbjV2uTkIDT+392Qe+BPjifAjvUMF
kYHWiU4BWwggOyAA/u2Xz4ko///PqzKtU4LNJjragZ4nVr8+9i7b+a4qzSHpjhkB
GIaSgXNMs1/3gbiqJSw5dcjQH0EhQCBg/5SK8TpNa48PFg+cVeaePbyacwkEnlJT
i+up0dKwrBb6FwgnkYFqfCB0qYVRQ0gsHCF3j77YRq3Ocf/oqfIXd3z6HT1PNkQ5
KEdADL4oOFD3drdYpNbvIApwRW1oxzGdYK6rEy4bBl15+KTJ/WtWW7mXdNfhF1oj
7mIgqKSDuQKlzhxVEPJWuHElpMtngrS+a0lLa/sD3XMhHbHRCUpwEUSeeicA6JdD
lnsJlBsEcFDUW7ZQUbHAjy7UAdQVpH/ugJExlTcalQ6jTHc5TkiUQJjCvHFT2xb7
A/M5m2ezMCZO7kj2Sm3TsAAsgDmbg0yO5apFZY2ofX8hki+sfSUkFiOeAaJfB4Dr
5bqIbTUubKUtF7/I9srfHvH1GksKn56RJPRcuTM9YXeqj5zBB4+DDOOJXNNg+vuy
rJ3VPdZv4A2cf88pvecsfLbqJ6yVOdX0ByAYGIIkquEGGQ0iKyBvvM4y/Y2T1MkM
KtJfMPl41V4XvYeif8zHxSUq2L4E3RQK1BhjBYy2seDA/zPXsmGL86FYd5ZiPI9A
+ImxXWKB13ehNg3AVsVWdg4Gd78CoxfmGvuvTuB9uwbLX7si0J++CnsMqXKPZupl
jgk4FbUNfC3ybNvRtBxVajPOpQBdbNX/8Pt7QoOtLYVjZmzNipX1juJ6vfh+wrOZ
BH8Inh+6REG5uxE+PwzY0FS4W1YewNucp2//xDmrbkHeY7pR+bp7Yi+IKmx3u/HN
GrNDxa7eoKqGbMT3hbSV20bzhgLFkUiUyMDKmPzrDKnVjdqexA1HxZSHAfureNKR
rslLJ4mRZ8JwWC84wDpdfhhMHzcrK8oU0prMZhjYj1JdDFyjJS9Oy/uuzUxDDOaV
gvimwTj//hITRHq/bi8DU9iB2tF3D+gShc/bW2WBqKfd35o3yQb43NS7sqasPEdF
ZQIqTD/t6f70cfdFTWtHQq8abE/Jive3jXmOeOu/xIF4xWao8zjOKJfHol3Stakt
kjOqHD3BwApkCeDPc3YgseO+yZibzjW5xk50VOGJpz5sEcuJTsCMtArnORXXI0BZ
yoOWDobF1HGVsvjdoM7IOS5eEiCXy4lCEeBWWRymOtgC9xEoelmPxc3mOFF50AO3
PvkclY1EvmV8WBwxnLEF4tx1jjikE2/MjbW19TlsJKdsexvZ4J16AMle+s/JoXeb
k9H7wlYGCLgNTDD5rE9FYpSSWRX/3XrdOYIOZ2vDtL9+6jELN2Xy2rkNeL6i/k0v
vDTm5nLGRvaEy4sjP/oexljeJHkxysp0gC81RApjstJUZYM+Bm2oqF34/22Yxx3k
ocktoORGfT9mCzGX+oy9xL9S4YiAlXF1ozvV84SmyPjD4WsLm+xRdrC0PPM9EXoj
BM1kns7wmzYy3ROlYrFkdlu3ardOzyKdGF4m4w/zHNra3Y2TqpMp+jjq6ZquoDHm
8gKKEESi4viPen/pcgwtPZgoVRPakd5HTsW8AMN0arTMQwWFx5R0lopYvSqvN6na
GFv4vHiqu2E4uSKncnj8wF84gEDvcjYv3k3WCEdKbghuRhE4unKhtWTOR2A5H94J
eTyPowU+NDINCV59CjIQTJeZ65X35yQRx87Wuxax31BU2qLkozewJdIx3MJiWFux
XR+eAz0DdNub4Pm6syiwIkvnyIJc9M/tkRrt6b/QaCA2SBWLOUFUCQ6dQopPyeds
jt8cOfgiiHj5amGeI1fzPgtehYXQSwBEsknaSVx/DUnSbYrLdDwpsbCpPPQjh71Z
obJgJGyzIYwHY9EDNIpbtSi2FoMFlhdt4Dxkx2nQfEgTNHa/UdWKRzmenGKJ9RFA
9BlUj3B6Mz6b8TdMWnoKRXX35zO6eK5ErXxcIlRY0Yu6MCMXg2a0oInmqPiFznoY
AVEWeIr453ZiixMiuEidCWDwtnYtENT49/lTBBRYoEMweERHFXPGLCAWAgWVE0u6
v8e/vQ5JxsFH/+EPm53Fa755hG1kVhOK7qNBd9eKm28Scb/Chww4KiXKg1+SR6e5
MI9AzX4a8Yu4S88Sb9s45/HmVXvu6AMY+/odNOvQ8w5ar2bWuWtrJs3eLeRXbr1+
mZj+w5rGq4mWQ+xrEwuZsWVXrKbV86iNfz/OyP6v9TRoUe+rlmwANiZb/XXq1tP5
CxlPx8oeQ1dfFU9ScwtuBpw0lq2RU2j1axtw9Iso+n3yEmg8N8MLJlR+jrx5YeKQ
/noOfevZ2g71dFCclJt5FaYTfJLoUJYPpRcS9Ru+3WyBWcwuu7+l5OzamuIOZaLL
KGMpyc7uoduS9OCDDrfRbS/8FydmqhYc+Ekh37oAN2UMXXddoHANlkAXncAcOxR/
J9olhQlJfujTU8zzdkwGV+DVzoTRjRNur4cqP5bUbwVODcVlWTL5Tp+FvvxCz+qD
7GArROX3KpP6+ss0xzq54c0GpYKlsWMDiIehoVTyl1mrYG7kFa4cnTJet1gr4HUr
BcWgT++v92vEVDG9iHW9FEM2goI8gNWNPHelCA63yG1P2Ok1ly/sP3ok/4lwcQLK
Dl8AyB5zhHrftzD23M3RvElOf3WgtEi7BzIn6m1oOxlmg2BgOZgst3Dd8TrPBVtS
u2jCXC54OhyzfPXoazXptGpa1IzZfcqRxP6wG4LsR3nAq3tzlGQ/hIKLppfjn1Mi
ghsvAM6sWQiy3xWrQXHyULx7122lEevtSiQ7LP8C+a2Q3ZeMMVNkNhAcup7L270H
rZt3+si2sJtzeEVs+HIE5OsrLRLSKkAgECbhUD1Wh7SDcOYWs64TVEkfAWf6coCS
ABMQhsd4DAUQQ0YvFJef+eYFJX2+bTfbYcGFto63X6GcPQlhmY7fIOcNkFXUsI/Z
JcRPTLt/31ms4zzwQ8MpKgZVe3NdB1lY5200oW4gTve23kfx1Emg7lwxSip/U/mn
8G9AOece6KVgYrdyfa3BA8QVI35TSqoJGNIp5tp4VhG1H2haViqTxSD9iE+0CKaW
DWIPgLgXHFDX7Rq8mGTzuOo0uV5+PaW9pqPWnr/+NwmjS5YBkaxiaGuSzofJFx4P
vYbnw7aGbuxK8IRoS0gKV8EkhnlhNLlzvGPD4ENXscKlfjKVCXMIf3irIHzc7CuM
iRHhlrDAHSACuoqKdxcRqHf9dlK3Loy3/WH2hJKIJTkHNrJBtktdDP5scCj5rdNf
7Fmr6f4EX27N4eyycbsuG/h6H6pg8vc3GqZ0qu0V72X6mYrTt6p7njUC7I/71ktA
VbPgBo2az2zciXdasCJUxXEKbWmm8Hmv+fC4tTevq1XulzHA1cTe99GlGOm0M4De
61W5DPSoNthTbNJICwx9rTaEI5rMjOTssRy/f8sp2yRN7bnK4rprFuFgxCu1W9g2
sDTZssj45UCCMP6R2XMLbJcMDA3yaX6RJM9PwtfPZnUCJ2o1dLROV1krZFXePS1U
gUQzALpMR3VKsAV0nRNlqcNib5JBp5i4EwRPjptPK9YCIRUSDd8wgcZu10lx95PF
f3O4bn24WZgRp4OZFH8f/11CjyTwRA29lP5xPDk7ISiqSXaCAcwU5Yg/k/I8D+fN
+LtuvQOh52jo4+RwQ5ylexHWC3OB1ySuPNoc2Gh/vOhqs0Key0wEWlV/5L62f3Y2
2D8PhgWA1yB5Uh2+NNASh80/nhP6B51nDUoGEhw6zRiuKC6/AxOWOWw8Zs0udhGy
de841SFQZIaPdGGw91qaol8SzZ017NIYHSYdg0RHIsxhgsAoh89dJHtOQf+4ka+A
tZNNG3zTA83enS1zEJphpvhFjN0FYLI21hNJfFXGcY0pcVAo4VohUo8IqVVnNMVX
0EexB12Lj+lCFosW8eFdMq4CuJq8Fa6HkbDZvX/FooCSfULBGs2loklPphOrLJq9
7nhVMMbr4/FvNrLEXSJbebPCa0/BbOx/AvXbkwROO6dFajDMEgqna1dQwWKdaShh
/4U7Q3CsYAjXqB4TZulbyNyEaHq4OWFNWWKIQWLKwOhAwSkPXDWPJxyAXgIFAhzT
mR85EafPWLEKrmuZIr9x0U4nAPVM9qsBj1+0BsJnUY38ee1eCiNeG+vKgV0nK08Y
1faJIsK3zfOY9QzONN9whX9VIBVlZoIH4P+uHi+NJiuZB5qSNU7GKDzaHnTpcdSV
EJTb9tR6F0DsDJSkhUbbgulPVXzyrwUZnDlsz+GvW12fzqFEFgGuEALnGkXFOTIL
jPnRbDOUIafWYkLpT+HPXBxGU6NCv11cG9vknh1K0WjxALFw6G5lzoUCtgr93X2C
hHR0GcuvSOTgBtySNBovi4RasaDson8whavCeCVqPG0AvuRedAZ61Dsq1CVU+5Eb
AGF36r2utMebJv8Zl/YpfaME1giMY4MlckDxyZftyF35YWoj65gnFZk9CWYR2KFU
WgE9Z3fX1gdGABUr/5lTJF6dNhDfcvMCS9noNqmUEI02tR8FJHAGAU3dNr7sU9K2
/BCJYgmBQUxrL570XJpdsT8q9itdVtsZqH4uBxEhdONeJAR7g9zsND+hPzZU06LL
68MbH4xP8k34MgiRIHEHM8zo4OCJiAtIrkhL5bbCSUF62A3QLVa/eYA/ZlPUCzQH
Vj4NeekyeuJsBY3l4TvWA3SH/2P2TN8ImbLkgPX5HjAG1zSODTZDMul4tmpgrI87
vMeANm5WD3zVPuKQUxQ9+Cv64UCtFX0BngAoeZCq8zW7uQ4XQvf74Ckgp6GsolSE
ZpSJeBmfAhn9OHBzBVk9+8qOJGQDVzrSWJdxa5gpNTDj6fOxOKLkyBAUmGSvaX+w
tphVK90hSx59jIcF+NYD9NSSpgfspJrJ//IynA7EuWXI2jvs64C534l0Z/Kh3qV7
7xczLR2k22cgWfD94zabbKpjYlbDF6A7k/JVFN67F0Z4g1KL+qDsQyKrXpt46gHZ
z8xdWD+4v4c2b7rVVt3nQFz4zXwyL7vuAb62CPY4kYdicI6kGdohPyoeVzR0SYZa
vAMTW7Bvz1frtsPW0Z+E8ZLjcQIE10MvE0dLmL3QpO+5wsyaRNWkuzMQkiPPLNh6
PJ2LCKNa5nduzWEYQiim5anFnSgT+DUCxD7DmSP/LbBsvvxBGJpkyls65xjorc2z
obVjsOxe8WWxkMXCO3NjxkUZu61O0cfwn7/fgyU5KRVP2Lz20Av8J20PUKaYq7/q
+eQBnPV1vaj7XKhI96ubn/7CZIrJo7YBpU5uLsKYExSxGxJqzp0X3Lpq+Q9azgVb
iXSJQwk4OaMtm/rlhCtKLaNG8dTLk78nUsKfhOA0Qzm5h4PKlku3iYHG7its+8+p
ReVyivcqbH0LpDmOhXul4bDndZRKYogJDYwL8MpO264X1/7UpQzKc2m5B1gztlAV
XBKIa4d0wx5NDCjDieA/NlT6zyXDZ8MLe+vcXvKu9aYyxwFY1Zm7HmuIc9JD9LNZ
38MsENvGYxdX8bxethUixXOmaC/kfeg9ZqE7KClDGyrb3ruUYY0914zxtNB8/P/L
tW3qBAmhP2I26QTkSn3mfq4HmUBCq4zESXduKjSDI79bz7a73ldh/vKuJOggbuww
6jDPIV3O0kkKRNJnrlzrqX8JYr/J1Nf+weehW670wLR6Bhq5/C9r18R7PQP9fWI2
3tJgBPE6n/UlfaKHTrr+SlpefbcojnCrFV9TSBrAL5EteGyWd8fBeeyxr7qBENsj
g+WPQ1CofvRkRzDVedoWxzKDb0K2AfhygTjOXManH4l3la9FkSLuikpaBSjEBuzK
YcJQJdAeZiJ342kLHkJOE5W9IiFeWKlKLFcNyMnOQsA=
`protect END_PROTECTED
