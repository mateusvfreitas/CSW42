`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
03jwQ1o4t8iD5NFhsoFAQYnAUbsJk1kr/O9Mbk7qGb0qrPfeOq4izSFq1stjUwoU
xVbpTrMKDttW2Ozfyd8tOhWp0j8NDnmGDpCJmwMRBx1jLlNyfvyKbA+A7/3Ybqph
EV+RYFM0crWr7jdLuG/8n/WgMac2RjLdsNgMpc6hizOdvmbEJPkYh+75sOnis7U5
qgXS2LVNczYTEu+DR9mBW3Go+m9Zqo7sSc51D37LOjyTRSA3a6ZONCLMw/bfaFD0
aHYpkw5URaKZW9Ey4y9rEItKx5siTeork30kPJX/pJMsrnEpAMKQHr5hyEgcJzzC
DNeRAL+CSoyiethwS/QbzigHAgMDRGgMXfZ/TGid7oGsJ3eav00nE7yzDsLGvb23
08kPGQhNBXBNRMJhOSoqm6325yg1abBRYjJuMlL+scHgenq80mJkJ02Lb+7wuDjk
JP2MuECyinFtY4J/LsP8c2dUqtnNqDvqfJD9WluzJzqJ2UUGzl/I6oPRhom/R78k
mab4k+2djGnADWRps91PgqqPba3YHNum3SC2/qHlUmiCYDsPKNfKw03xb8CTopKF
9ZpmqfFnBye0k8PMxQcZyVox5nRnHb0p+leJxMSKUasSGEhGUN0vCuyMzMIE0znw
waFf0E5q6tvOdq/3phJr/aJK2zDpLLeVMR2K6fF37vCg2pwJe+2yL82i1tL0c19j
nOpcWz37kiXwmkUIanChdyg8w7jsyfSK4bmx3grPOfC2Dt233K72EyS5h96s6ADX
JvUvK4+UIhGikIc0qRzdLxknc+eKzVE4DWkRj56vrffeR01k5YO74iuppM7ZipLz
obBrtffICYTnN89C+60pFIpngrGSzw5fipiBOmpAdOcPn40siZXSPXU+/iZEsHbN
boz46/U2D88QswICR+2fCvNZvvHI88tFLy6DOVgDPqfyLpRD4GLdndTid6BgsdNo
DMEcjmIf0YwuVn2FBYw/unJQ4a/1SCo28SP/6+ka7OMWXht7Pe8v0NhDrfw5CFca
IpOadwf5bE9SRQzBtYvgXv+80T97JiUlUr8BANqhUkuPds1pK+76p4H9DwY67Lo7
bBvn7YhXqfSeTzB6trrFVXS+E3nL6UFI0UI1h4wlSFzdDye1VuR9SBD45mVTYpfr
oyEqaUy4+XFAaxRfGvKg2pPjOFSirCtcdEi33pxN/1aeaIXoc0XlbEMMZMMf6mI7
BVG/iQ5+EGal8T6RIejtFHpvGMxUXl5UpBfXThfP0JbcSYFbHjjpfBUknB+ALLmx
wbTGEEdc6YU8wSfti6Sdl4XvzY+d080gyKyIvwe3W80ITJi/6B4kSqTyK+Hss4m6
3FRnBJW1GRddszJ7Q/hMQ3GybSW/PJ/9sl3E8jZxTk+++v+JKCQa4d21Q8eyjsLg
a5mUWN5U4p/JtQtIMJ4jAZ5lOGjYk6fMlj4p/jOxMEbt3F3TAARUchz2pbiBlMy1
pGLF3ZP7ndy2BwV3k47b7Mr/OnLEcbgEmAhYAUadmYLCJC8vVY/es/7tevJyQbiq
m4hMRczBRuFPaIaVPA9eomsqUkdo2S4NTugCgaESxN9G9aLzTbeVNrAggeLYAncZ
ke6z5W0YJyoYshI+DbVR6HlxemaSVdGCpz7evFjQJp4T1v08SLJgYfxddeknOt+V
GmecMUE+yliQ4iQDOz0rw8V+OUVJIHmTVTG9ustDr0cv0Gh/bX6JPGNIHYceoVxB
AtmxF1cjqTuVO0eKnq/v2WqkSakzTMhSXkyM+UEnbw8A0y8oPII4K3YTkjo6Z2If
8n3JeXrQBaKNQmXBvf1YBML00PYU2W5mFR+poCYcrq5IB2qGeMp8hDrBj0zLCMEE
0JyWqQ8ItsXvAqf/wD9u7muX/mr4XJpa+3+UxhsWfwZLNaRUKhXZaQ3zavFHSTs5
OLJXJzUBdVHkRiTzHu/tNKTGRkldtc60Jtnc3mk4ABOk8c15lYRuZSqSdG9dh6hU
ATLyuMtmAc1bqP1qyrzKuY9iO7nrybXRD8IfFfLZvT0E9VrLhD6yVSA2nrsb/oAb
1IElZRuzkC8SGbwvTRbLqBAGHunXYeOOgCRqFo0BY3QNKTXY/H4LOfw7QRCUy+A+
ZYjw0z5gFlQjv8urNyccwVbezsuYTCv0F/6gZ22uSo+cHpVNLGsEXa0QrtbA4b9a
sg4T00sojwGriHl1ef/8cjpJ8hfO9Zlsk8pNhkbIxqmjSVnn/OYH7b1g1XCXivPT
AdM2v29mWQ9ic07vw5eu4A==
`protect END_PROTECTED
