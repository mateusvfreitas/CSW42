`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q+RyIjWKCkotbkpjnjLiUnSDwrsWOvzd/sOf8mVcnTzBjNfQ8f9761dFkFrdvIOZ
F13RfpuEiLKQGxHFoJ/4Mm6yGzzOmvKrP876dWR1uUqvzP1YdufNWl7Wzy4jCAl0
ysBhJCINxePXNz9PJUWZaqxfKb6Sa07ANYZp5850FBMiNiC17VYDiYXob7DsMKh1
RR4WxB7B8IV3AHattNBcZDrjDfaULhE7nDKihWwf5bS9j+lptNuIgWNfiTz+FU1K
uX6lS2zwXriY9E2PWhkVVOS6nlHIJic22KZfH7BtYh09ZG35jk46BIFTs/MwCNC6
Mdgngk8Jc9vpPL8sbC5DmUEsE8U0PtGeIz7jLen464kHRcy5Zfg8UNVfnZWW7w0X
c6/wAOKdJdw3V6bJ8oQNnOTjdnhCtpTbUq5lCPW8SHJLVgEZa3Jzfe1x6xe5d41S
JYmG1qbXPS5BMRLwNApQjxmF/VauOVLYL+zWxDVvZLJwgeVhlrRIIxZiIF5zu0aV
yBvFoJFEHihKm0Jx1LXJbnfFJmad2NpPdlc1qOjWWg6vmDWEaLnwW9/ZAfzqMB9V
8QSnOoT3SHtBb4SQsCk5xEYlC7ntOR/BHe8NYcQd0XKDyJiaHhLkVqHovnfwMBy9
u1N4+gXTDZoyc2gmR7E6G4GeK5NzxHAMgsx6K3EQJ7LBJNigxbQlqVEipZchx5yZ
I2W+/99ZcHKSAgoNdnAQZtEeL/1MwkHop8RINW2vZdBLvNmDN/YYOoJDD9Ih184F
/PBcQlVFH/uPzHRHb4ntOupwzLjR2hboPxBBIzYOeGcJu7KWA1S4GNd/EiiZSPmQ
bzjy+fFKwYXPlezLYB/6T8y2TlzzFHDF3sa74wgKHU+Ki3Z0XEDAVJNO6vwf0KjJ
q/HawpfIpql6PcZzvznxWuz6YXdEKwy4zv43fIrCYKTxpvvt7BQ2gWFeYhxEOdbD
dOF62EJfrFVUkwHggbN7u0HWeH12Z2AHaa07Y0yApn94UXTT0VCOu6UIsAj81cw+
jsaG0ITaeLkJUTLYEl524TEWRRzTy4WOGVEBuoAt/KGkznQtf544bcE5BrJOATYK
vM39sj5iplJ8gRFoUHA7QlinAYgk4WkjVIaI8SNG8gsmgTdERXd2Z6LtPiFQ+m6D
WonzOqG41LlWyT/6pqFNmEc7hAGGpRl/CYY2Qw4nKbcxY4objKGtuR7BDfQQSSO1
hX6+ReGyGQKYJvUZIUsrNAvkC8JgOreQYbMLRkZi7zL8jJwbW6eSTSHJQuBJFWyo
9w5YpyPy/EqRHGWBfHqXMnf7vx881WbHAvDjIKci9lXBt8lS0WraTH2KcliXWvmu
nlMF2EY5oq1BEdHlSuaLF9hDC7VDTI547er0RytQ1zCDdkI3A1Tzw9isUn70ufkP
NJXnxVsYN/NbPWPAAVcNO8O+FC1RdQ474ItnDSV24ezLsqSQkvdDcs4rbN7uMCrF
XsMkSB7fl4GKblkn36ngHuwHd9vxyA33bL7NduS+7PqQH+hOi1lT5oFrDjWFGKHs
DTEfDIRuEjVKHV/S/lGSGuFl/xCSOIbEo4LxJy0ISAW4KL9i/bWR1yYVGBkrjW/o
axkK4+7CrePeXNIEoNKZ55Z4DbpYS76Y1RNN8JKIopvHihFt01LXfgnJpPXZpYYo
X+Ncd9XNpZLRGqRQu9VBJ/BgzAFxvoKOK8HTAx+QwJmZv8jS/4IFeG6AYR5tMm65
7Pn3pOTvOtrPc1osXmdVZ4Qk/943C3pfp+B84F86QURDCdOy/D6Vr1CTGEpa+Bn9
fwFqA+u4nRuCv58ZpUSzkNcyPGttR4372n2CfuRSmrghGZmibWAAaKHYAMPeMXjv
e1FzuWO0RIrekF/tqQ1KKE7ZxN7RLdsOtvILkxeuutPTiyJiQkUMPKZ6qtI8UpCw
Kjs2pzXeYOXxt5ZsVn/u4hFDclQeiA9eYegfMuZcA5EW2p6JELxWIJ+7ONNQ+G5D
R/U4j9I3fBkXFWEcmFI3G50m5dG4vS7VxytHYe02+crABZX0WVlG0wKVJucgEW0p
pHjiMPreTKKIBDcjOKUUyGJj9RG/sGwDLlm4FAJL6RtP0Ihnzjv2to4yY7msZAcW
+N+N6RDhIidQGekUPa5Jiy+tidgAyKLFZCwKdsAGbG738sJIi0CTnPbgQyu91wqy
cephmX5R1oJKj21UykR5D+THwkExw3882o2t0g0PHT3JHmisC3BxXg0yPRqwXF8w
q3OEtRkt4rNCtwgo4ZL/o30FkIDKDsiRduRCKyOq4HFq7GyGrNaIu+FKsHRjTwON
DVM10GjaDdKa4nuWZKChQ1iC2aJxkup2VZr70MYuDgd4Rz2t0HiMk8vAPNUOk4Vo
F/4+iSdATmlrgnjwMNcmDT7ledqc+veQzl2Dto/kEjxDv+93pOdVGhffJL6t8mmE
fckVuSxEa56fbTp5NjNwsb0qNwcOXqJBO6VeVum009AjruWP6c+r5/viDw6wUr/g
WmuzDIF7NyIf2BYZTwTzPHmkkaIpR5sPPFtJrSF89beBnqlrn2kI+V0U8Oo/INIC
+Z/4GNEMJ2XjH/p3QCFjplwXukJs3a0hdSZ1e/ycb8h4VRynVMBRkcV5zc70lnkQ
q2L+eUCJC8bOsz8uO58fRsmzmseiX86FU63LncbERrV3e05PZfnuM9sItZWs8UsF
6YgKLA1eyTpfDpRvgLDtFwLILNZTesxfPLHo6bONs4K0SsC5NGKwrNTB5f69Rone
VIkVuuTqfo/F8JEkA3STWLyNrSEwRCddFwSMQ9YX3IFw7qSz652/fJGv7MNF0MId
ejHpJN1xXC3cWeVhmNG9+9m4eWNlnX4wUzK6qT2U6iiQiJ0RD2u6+vvV2fbHReM9
nXZ+mxdMrSoRUdQ1HxR2631v8OHQBQ14lgJdnpvyYXwBEQR7ptHI6ojJPt9IAHha
RNS569/qYWgtuSvHZHn5cTMI/Dl+uxHtuBiRUd7zBw3gZjqVT4XteYQJS6rKDfmD
zkxpVidY1MdQNfbua8CPwZegeH19XKqDspdOrYViwR6bOvwSMLfgdG0jRWEW8Qrx
RyVU0XGr4wzifjH/mNoRxRS7Jqnb5SrohKEgjWGEkN39FARVOi+kTHWS/Qb8BuUV
+HjWlgSp7/KCJDCVizAisxDxYDqAU59ZxchFNUfzzABKVp0IoGuCt3zKK+Jeu8L5
ZM5MZoQTqHOuse7okablJxFKwgUD3JKUUU1u+Q8beG1sr7MawELyCYDdlFiXOUf3
kcS7AZappmGP304rkaVphBt+0CMBzibrMkcvWw8SAvhKFrmpY/i29y85va0pI8E+
aZJHiJRgUoQL7okzMZJ8gOWvkGpuibhu8VB/iDAsmtYJiMH0AKGkT5EH+Qs9W0fZ
sdzqQ6OnU2yMCqA8YLzjB4c2ZeHMRWpWbdd2v8lVL4oi4U9skTOA0EMBFtU6k/sf
AA9Ldm7Siw82YNtSWUB6FjHGjmKW1gUBXUSree0RJyOxxxMmqW4KCoLjgBwbdPq8
pWwXL3sKDr1i2FhfRaqZD2DBc1LIk+nBkb2BT62hvuVwwcusN6m8OPaOaLk0jyhG
8jLw7CBt8Ku/F3j2VMuExMxfbC5UbuwUs9G9z6ZzedYoFrgvl5f3wMdwqVCGfBFL
3OEQhWLmExkbgFWN9rSqK+lITgAEO8GImUCxoIbFw6t8hml6niMd2t1PDZlXP95b
imEvH+up0DAhUTnRwkkJtT9plbfCKxrXu+ZY5sxzXcs1aF5dY0WYTX3oxzxLH0iH
2y2yTRU5KWytCZ2ZD5oaq6HgauIxgD7jrJNPe5fIszNHnDUal9qQiLIeXPOj88EI
/4O0e19ZBPSreQxUb3cVvQqrTNDgkaBAkLHJgAmXdhBwbJE7j+ehJe8yHQKmXesZ
eSTAwwdLHXv+spwj1/9DbvyoXnRqfAk6jEqcGdM/GkVkC1IkeISZSK6adU7wZtrK
n+CJ8mFOBwF+yqMaV6E/sxr5BB8VB+H+ipcuBQ0C5kSkUJzoO6MxTlsQMZca7yI6
OrEWwrlaGEybAK3DJfbesYmos93UnpdWj6H276CU3t2OM9D3hHbGKCbH/VihCdhI
pEDnbZ2AQif8MYQcNlND73ko9vvEsOZ13tykG/KP7iM+Qb/VSqG3kXpnVnzJNSnw
axsVbNeTPWWLeQytAVAU/aUu0WeR28B0hmXXaBsF1c8kNU17mnVdk0Yfa7pIqfP8
rLlxpC9D8sHaGvvi1b/1D16P4wzKVDOyFYGFQiNT2mXWFK57OrfOXEDP+3dYdlIv
1RJQkTNlMl1f6+HZDrYMhB5pdaYzlmLWnJYNq1gMIPm3sUL8nAHS9qckvhYDx5wF
6vCLIAF1MEDZgWVXlWNGBdO26WJu0/l58komNiYK2Sktgf7KKOAueewRTBYVmXNI
f1ads75QCWRzU4rrVILkbpwcbnn3HzfZQRVee8NcsHNk551ZQ0whTbsREKr9/jSM
xMkpaHG0U4FNNdxVID2f/683P44CcLPY+pZa43o6k/UH5TTgJUDEaEoTtv43NqnQ
8KIo51JEPJ8k4qQO2ZIw+ZnH0fOWWEqxlvAAidVxj7TAS1IUn3oklEP/6f4z5RY8
CpjQ0U1zrbIYtk7QreKXkHwl/iRk6LiFoB1qPvgXChV+cClVbdCD8/NrhA6eTiKk
p2bULSP1DbW5gr+jUzAIGxsuebg8FczEYgUQpQBpCqYvOEspRwgJvPxg4cPJiLgr
UmHoXUTQWmnpH5NOvx8hXKwD1SKYYAwnNI+f+aJxkIE+shUjWPTDu1SHi6RF+MTk
iwzNzxyacqkO3Bjf6AqR6a8/SSF2Q3NucV5/4u4GGvTbFeE4Xsvt+CxbCKBe/g68
ezcS3tZCgfUBA9b68HKzBjFuJtl91sdV2uCpxoBX8N3yrUETXnVi4SoPUNLhOINn
L1rtcVVIGeEF+zJw5NKW4pxvZkKcyPoWduT3DmbNNnXy49RnrMkg12dyzj335JZA
ORZ3FTmNmo7643faN3n8AhLVS/IcEPTb0nALk+7qe2PZWTAhVHxVBHsCYWCeQ9i4
gc0ANYsZ1zpyCtEG1SagvfdBcwE+SlFn0Xc18GQD2Q8J/q4IFMF4lJ81g3XgRNNo
s0SAcCKtG0mGANH2o9qHd0xtChws/4Qt9viQiCddIMOjDjCYLV+Q24CTahFkNPIY
xVwZIUjaa7iim/2trZ8j9g7avESPufjddVzSc2SFR6Vy5hYZ6Y1dodQ1esztP4EK
gAeet8FXQaNlADZPS+W1cZOHDF18J0I1iDnZBEpqlkaTPfyuxVVlafE7apAkA101
wHMLhO5zqrwKIw+OqfzCleVq/1l+0zO6FtEBJrJsw89ai7b0KS6shYOwkEnZDHNd
FYNTZ1JHqrf0xA+B0oRyNgoWXlXGyxwBu1yAmY7FeM2NBIgKyBTn/yTEoHn7TYhU
uLzwTZ/OlfK50F5uL4e8ZVByv+tKjvxSHRCWWZu+nSO/pulQUhlKNJeKmgvKjmQM
r7WLfYg38goJl5+C8zWkGP8u84hjGkpJh0rTBFEfr6HkA8f+hlgtYWE/JpL2WThj
4dNvQpd1XvTWkfg4PTnf7VYEc9riOEqk4uOJrCYfEuh1fEgie2z4QjK4QbdPQYKU
5Q+p2wddwSSmvnr5zLtJ0CwEEnggtHIUgKspm9sLlxk8CXbZdL/Yl1mmfZRDx/1Z
YLwlUkDTtt3tMHU4+6mIuhJ7P6dLocMZ2pM9grzp3J3+cOjc1UvfQcabGkWBlh0c
mkxfI4Pzfc7Rt3WPqshTwBjKLdacEzyRQgxG8FDmEOBMS9JmeitPutRfzSRbyELF
igw8fmZkVMyW6gU/qilROgo/Jhxpts5y4HvJtD3aJsYfI1gHaESCA4sD4TEXBDW9
YTYAAplBJ8XOrrmkcOAaSBqVRMBn+ChQkSHpl9H1oDv3cmORrw2mAEUkFSpPMsB6
u/O6155uR1gV7ZDNo1vyClAstaw8joOH4xySm7xFTprpG55KiMgK3RRjo1T1x4r2
LFibUPrWp7VcfXTa5Xz9Y0O1WA7B7Dhbnon5V1biq2hzajT1fmrYpOJyG6JW9JR0
WyMx310gsPlDzKGjf/XVzmYy4hc8KuMbzeolUrA0O2wt6gWTmVbI7kS6r0/ZAv3B
kFJcHubH2FjfyOGsnheX/PnVpU9gr4A9GyjGpNFBSCLxZ9SRaIi1DSwz3k7vlyo/
Hnhf3hDTaeeqhyAnVtyQe4+p5RVm3qhzJ1P/ikJgMxsYqE8XQheGZmU0cKI/xLXe
tslPJ/bRnYYwuJ+pEo76U4zG6+iBKAmPSz+P80n2hacKMtGPMO9z0tMm4489aS8S
8sWfbkhEJL6SWFT0RWY5UIN1BSadnrrqOhQAjS7rMuDMr/C/ReMTpHLpTr9MJZBg
A5NQvnYNPu5NF7pj6IuyoHJ5FBMTiIDJ/3yy0MM786v+iQkENyCvsbYRt62gK64o
rgG0vlwG4hX4vYvPhEZUblQ/FZf0ZWSOLjv2JnuZBL/AosWqiC68RfeqClZATg4Q
NX/IdE0ankMMMQibeBTxzdqvZ/bajs4JhARaTLsyS38QQdz5duysaogVz56ptaUx
x9c/93sVA4rbrAb/VyJE/o0E5ln0qTiO6+r6nLnIS2JVryPgYOM/9ut7AGbgVxF2
Z86EntsKbpS1BrAKLoyk0W7cArG/EdIVOkY51fCuzUc0rpiaMaaJg28eTTCmUNaP
+CbWEuHka5SICnlF1v/W2dhq42MjQeE3O5s74F7TZfXssWhJAB7khj+YChMzFBNh
kc2xWN8H+ZIJCLf0czsdWHcVGwU4LKY52+4f04mDoUG/0Sst9HFnfMeQcskQkpva
DhgmSWB/38WS9DlTKIDLBmJQQJjrUI9PUK6tMqfFnI3MU3RUxxY8iSONm2E5kJSH
hFkHPjuzGY5Cf6VGJ5Xs7oYh7bOxAb4/3SJpxIDCl/SMqWmmY4d14hnufPA1mKxj
7FZ92G8X3U0s13tvcQFKJWVXEc3CARVmHmpBuKM4Ri4FgHQnNUxaQfeqHwFrYbQE
pUc6OmXw2LHvdAkz5HvT4aCs9Tw9khbzIu0AyyNUWlwPV4DpksEg2k8zXRp7wydZ
Urr66Gxkj3/kYEkvBKMArt+NX0EfFNGiUT+pZr4SdjXQFHhmtJ72GMWs2o29UA36
Er+chFHPNWLMf9plJUTeIASUWCnE3m434Wl5tQgpretO6Rvo5a6IDJ2Dh7MhsmtR
XhgFmP/MTczU/WXmdqs0+3UZcqhA6eonOx8Xzc1X9Pm5cYrso2/uxYhw6obkaFUH
2vfWqwKkSczE0G1i37SMUUJAwK6neUs1UYOBWq3tHPpDRU0AM3CTkE2uVuL890Qk
D7SfcEzy0R7y6di7WGEHDFXcK/rn6RSMX8j8XjpiqJa2fOuG2SSj4ipH/qaMeidY
pdBAM1bmi9wHl4S6aOeykZ2mSB7oijXGtEUEsTsq9w1jawZ+Qo//6ejqb8FK6eZV
nEUJEWu8MCOUEyDh80a4ui2rRKnyxcNNaj1XkU4+LBbd/ql9VaFb//YX7eipOzl/
Dd/97JE36qWBTtG4cS8CKpKxzubqRMkm0fjYvct+LK2etkToeTqPTEYmlWZbOAaG
oVHkiTR8yAVjepPtJBLLKOdZ8DOH+/eA0+a59oFRfoUGCVb806w9oTuIV2LEUPDb
4SKHA0KUImJXjHIsOxur0tiMX7wLuzbYlmNlRWVVqxCxuleZuurd/a1iclu1oCWA
yZkv3mhLs2IM7KGTcjSELYG/OzDzYaOZoPCAysr4kCaBKuAnpDCgnlJt9PZwxOR9
a+vGgb3GvSuRiqu9Y1oEbCalXunJ2iTUUCUbTGWLdZ9S1zlQmzXzNSJ65q5rKxsl
DT8B2gD8Cqtd8/eLvEk3JzBKF47S0XgTTWJ5J5jHRJFYsGHXLmUTAyUBJEdIJDif
r7Kr8gawHh1RmbUC4FpDen5GNQvoDTS/D+Q4H1TU1ux8I3otk7T5wUtS5dhFx9SJ
cB/Dl8xtKSk9X1VFMWxeezpLoAjApd1F2riesNlieQI0wCMJlLRUW8QWg8hxY2yr
6f35ccNNhaMDpQopNmfdr9Atqcf/xiIP5CLIcilcY9pd0tlX51R+gjAX+qq7mtaS
2U9K6KKxWfxariHWo7sk8DgFl4f6FeoxWHYkW/A14lTfKpzgR1dKFMDaDsnAotee
CosVLq5s8YD7GHLhXpTUNHTc8MXKxtEEgRpT69om8q+mAb2nbag3a3pKBQkGEiQB
A6THMPKYyrFyY/PP3+2j9NjyrpMVJACKJSODhWJs8eg3sa+8m67BA3LWcJ7uYg99
1xEsQU5X075VJjV7jha00k53qhYlPYdTTScOilRI2ursnfcWDbobXRC3I96dgRWV
bZXieZ/xndmjz7uBy4GHhAIzNjqKbcx1KQ5h4BuDjTal/bixSHinmmq1mlf8TEjR
5F0EylQbBtdc3cDe0TXpU420MLvr8VDFFeMeo9xu8xGQ8lXkrS3FUotCHUQWwTRT
hz/EIhYZkYcflNy/pVSMPlRbGr8I1+AXLiMu82c/YDhuJXBGrdDlX9jrQi15/VhJ
4aYPV3w/OJhRDPlb2XgJJfkMfozDRCGqsTkYqQfkgN5391BE8i/qs9wDznn2Zgd7
DymK97yM2j+AN4cIhcn5ebKLN1FO362z+iUJamUKf6Sjn7/9W0Tx0mCb9MFy294y
YCz8VV9QDypXtTHKjPMH+cIBCOMotiCEEg8uyxKdtdnTs9jY5534H4mJJhRhe2v0
0JxkzWmVseKaFhh4mpngWFRzvDifECb4UieT5AW8qYq+Ai6O7vccy4uN1oLeH/DB
4Mk0XvR+Cw9h5l4G35oVlUd8BK2FQxs9v11sQY8zeTZVhcyGCXVbqZ9VmRNJ8fZJ
T/AFDIuaC7f1VFqeAz6bxskVg+fYM1zAoqO1jEpm7oo=
`protect END_PROTECTED
