`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
WEm0KnD1VOjwwYwT0/Eontl67gkYfnB7hZ4BOhlCMND/bfELXTci0xv7dNl2lock
NjeQwJv7H+/00jyCryqbbf2JfifwRDmgnPYGVnsTEFOv1bgFIv92ZpOoSRzs3BS1
Sctru5U1tY0IgsX1XLJq4rc+3Skt42HCMEnO2GGqYc1ThRk+rIoosPh5SDLl0aif
efeRjWk9sLFLOjJMgF3IXdnB6G+rThPYwf0/3q0FLi13BDFs1UDgYKqHcbusN6iY
7uONdiDfQPSYGQTNSwdqilNZB05anHkmIjF7ZIDieZepabo/bIeleFkqAQ2gN9lI
pAko1QmGyTZm6i+dz4ytdfVVhZRAqUacg/2WuYic1WEon8b2I0dJPSoJkVz2Q7rY
VXnlJfLVeoDD7GzkmgUDPy77/KC+yncLr4t7GjlvkZjZy9Ks23j7ooJBmo1C2P9o
31wTHesIyVd6L0SQ9vDg90ox5OYrI2MDWkyznqg1D2YyTgR435otrtbvmIpVgSFZ
1Dfc50bSrxLmPfkAJQGE8FYDizw7i4Gj8++MvFuZbPNhV0mGVv9LDF0RxhWjhcS1
osUN6LyO9xwUYQPKwTS5PDjfDdkznclcZAx0uoKsLUg2sjGBMhY2+km8FUVg/RkS
k0Ht5RLI2EsqMAKXmFvuujlk1i0L48SIfRcJkQy4nL7wxpY60qgTIAx+3w/YEiiC
gLxaAQSmiaZP817vD+f6HIEiObXFNHm0goJKyeDN2yxgAPk924rS0tlTDdNbH2r4
51g3PmyXq2lD9yPvjGgrKfDJrskgAPGa3f4XKNHVHWxcvtLvu+h7POO9tz9wKibV
Wv60SI9T6J0/ZsULNpr2jZWtyS7meYowfD4/wBQ50TdqopEUqX2mBi0I4YD6bqCX
IWV4YEvPqXNH+SuBLKSIUH4kCb0mxVbhqqS4LZY9F0ZYG1Tog9uQmwI20DLXhsOV
BLgxq+xthd+S3OA1ZjcnoCCMqYjYisl1gqMcODnfhOwk+6fI+TZySkNMKiPLdZr8
pgkve2kewNQHTGCUBHjrjU3ZpGBQRiceSurOShFSZPGvmyWekX+KyGo5iC7R7EKb
3pWAzmefURCES7QXopaJKSUTMb788orYo2iJABbPwYlPNrIKs+9f8P+bkYILsKIP
yQCaa5zsAfsOdE2kN/adsqWQcrU/XTLLccWNeVv4p8/tUkfBsoDSl0poXf9d1ykU
pZCaOmuQtHONskNt3Kn0o8yUWG73FyEvgmaJ4WwnKqgy+t4oHfslS9WqjAGAafNh
BUxXN3xGYj/MVSYel/JvphYDVClz2JHAp+8T2Nx0Vr7jHajdOC0sP7lCiSDLacjf
s8EyKqgh9Ld24hRf0M7HOkaV1rkprWoK1XVlkZfeR5rpqLSgJAQPVN9u15M/2deS
vCL0ZXoUpIyFajt9j4N27hJglFjp6UWvB0TkbZbKrIqtFewp8q5zjZYU3VKoHeSd
U9naGRcFNnLtR6y9YhoMX0hWfp/736GxIw9guxAXfW29embJqDC0wXv4whdXx3VG
IrO2NNxNDnHPG2xPlFbNHZV25kk6C53fmjdPbcsbVMUSvfcIYikhcbo3qgB0NQLx
loWVdyluHnmFXgEG+Yt0tG5a8BM+cWSqgcjT9xmnfmjtfqBxr9yG48VjYkYwcjzz
CbTk/AoUv8CkzHTyutBW5Q6i0bj8lRmL79hLzkN1vUN9EcQMhBs+cQpffJrOek5X
m6dxCuyUMKM1CtlRANt0I1dNtPj+fPlKK+VwzLef5P8kv5PgrM+Ruw+H3uCSeXoH
x5i6XnQk9VGI05aZHtog/KusRs7erZmpx3olqY1btQjSJqUovIYXMAJTuiqJvWB7
3RxDnJgLoGkp/+aTYkzGwkpzkbWvX3OYHcX3bJm6EBOP5El5DL8Y2MvE8732tn2G
GUB9OQ4D8NJMiWo1bWghbGVYZ7uVo4z11f/8LIEgVxeNsvoeWROwPz5l/ZPlkSFR
xMe4HgU1eJwm6rDrst378HtonH65cdHz+RReMHvKJ05Xm0mUN+Wr6VwVgi08yfFI
`protect END_PROTECTED
