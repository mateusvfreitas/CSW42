`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ccCrjsuyGjqY3vqnU7sWEBsJyjZzaQppd/yR5PUGHNAv+zeIq7Xp6JgkmaXgI4Fu
iy7JP1pvnfCwvxWgkNAT4thyl585yQ27VA37Ed1Knr0uN2u0AyCjwOZzap3SbB4F
qs5ltrx0wV39FDFFFdP/tmONuO+AQp070fwQLFYgjtePHuZH58mMVunqQA2AeaNc
ib4hTXLC8jaE9ApRoCoO2LB5Mrq7uxyXruogHTCf5XZEAa8cIviD9mz2KcmUiBOv
BTWBYuxd7hYBX2Dhn0r5WoUs0AoP93iYjPzrIuwtZm0GptmEOWzYiWUuZ1ScwKnz
POHT/qnz2eqqH6iA0W5tH72OBiOiEnhyzWmWhUbm5BrFzfvHMMQ8z754ywsD9PMs
njKbXxn2mZG7WRigB85OLx/HowoywOAr+QJocWab5MSLxc+fZLPlvMaNP565eA2a
d8e64rjId2PPkat4Vj2HBAsz8DxAFrcmMMWIHf3mvynSJhffsxHqHUEQ6bNEuyih
sHnQjXFmypMJal4NR47wnnjcVbP8/w9KUjomPPUfEG8Jb9Jk0nuZSNAvpWBJdXpr
M5oBWPtlkItN0zKY0GwnFn92KCDhZS5hiy6ezXYHvSidVSuAD01bSxs1c5Fh4V+Z
8uCIKGYOu+QZber2NWeKAon79WwjA9obqr+VGTQ734woCoiV9n77/f5I56JayEcM
olMCFMzd0MRhtJQdMx0aJWqt9KsQu3AQXfHTF1fE7Ns=
`protect END_PROTECTED
