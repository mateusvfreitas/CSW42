`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwDzD3rCaPsH5oP9eu8FgYrlEaDQ6WuvmSz+zSKccma4fqVpBA8v0dB8ggKlMbcL
/Phm9EEiv171KKprQQiOu3ZDA3tpZIfb1jJw2fxJveFnlwsYUx+sYoxGq211SFKp
yYp8Rc+6C8DzKZrxBR5Q1FgA8v/qQH7ChhuiMmbexPKWvV5iNgwoPLvGNSqKcLKA
mKsXpfzKXnbNcLZKMAQItt+LLl14+Loy+EwrFW1oeE7HWEinXAUBIElFeIGNVxAn
lsxKOnjUjy67B75UHnBghXhxtjovmPqAIQQ4Aj9CQoXA4A82+QrWhAwuzHNL1wdj
UV6OGicKtBtxvTh9luC5D42kTPTuHay9PcZNhJVP1IYfuNvIvXL5pOFt9Q0pB0E8
nMQhtiqoWjAAiHwTqVZT2wBbsf//4XIdzRRB9cIOu8wfIacidqX8ArVYPsQGqY1v
RQbCgOffXcxDv9gsQMtmhccbetiWTKoEUzLKoWc5sxPozsIgUzCJTX5sreQeRuGe
h2zC/cXyJimGRjPMlM08RHunRGLNv9aQo+6Hm6EP5hLsd2kaSPb/CvPclCPSANIv
T8bveKDXTK8u7SnUsYA+WPkBeSyNptXQL48gaMipqgevuizvz41bC68/g01fW+hd
E5vUJ1zuEwplfMb0pHwKJrd6SlLLnMt0igVrsluGVzDaaZX9BxbOoh1OSgOYXJQ+
iEp5UoGVndD36pOho/aSGM/0u043aniAQCblbdKbysgR0+MxLNskwwYfeSAq6uEy
KshYBB2DjqSV2tmKq1EQ22FoFqpz5duLUea6dCZzFA3C/YmPJdGja1sE848MCkgU
4rnoWk3gk3t7WO9DgGKx1nQchrhe+CbFftCIAooigYMsGCBQISx4FeNmKnRFxxLH
St26QFpLSLTtSX949bH41xIzVz8uA8cqGx8swWbhkhXdoh1aCuoYpj3FFDKPvKzB
ZhnolrGPgX3g6Syh7vtZi2QECqGzNQ6J9hw4yMglIOarjBg9Zr9Q9hgLSY4EXzv9
znJeNo6o5mtPVCfsCyMPxXdpgtYOiwtQLKrw4FBpzADDU+QFOwBNHkl9/YnMFvfo
W0nEEwZL9bG8wHxaM3Xx2DVz1j2YbGihmwLPHNBcdfStNaW1SuywmAZY8eCASz/b
LG/Er3RQ2WgofthlYFsW4jkMElhw2VxRH8Ju/vyq4hwrWiCTuEo+UnxMY9LQajev
BfgzVBDYw1sC/fIBBOt7F4hLpbrS2ZP4SrGdVBnjDqogORb+d5PthgabQW2mcIc9
+VARR2lfOFTuYxADQsn9hx4kjof1uPh66uQ3IJLHleC9QQku3uzYQLE1RkM3oeDD
/YpNRahE/u6zo/xmNJc63eAovqckuLsffAXtz8PL8GyPSInujfazu5ctNCkOw+jM
PewjNXB1xfwTNOKVnsl8QwXZq8qS7g0ZiD6swEflNPCBHnKOjfktvOuOunqmdrql
EGO8Wbw8ziTU66cdDXn33K9q1hGGTBie7rXamQkdYfHdvCAdAX7egHj5SH0OZJHm
rtdTJ9ewD9lbK2Gnn1vtAK885I+wayrsmTKIdct/KpuuHPUsYVLreoJB2n7LTnJO
5i1dzUBPIpjxHZnHDyE4Ulx0SMTF55B543c/Qe2FcSWbUjD3uWYQf78NBTrf5m+1
U+6zDGIVcryurGAKm1NNWAKWtylbmY/7nlUXbjIlzm33wUKbuiMfYZO5xncK5Z90
y4MtN+zDLEhs6J9qTczTv4nW0Z/INz0Ok+e0e5tQJE/WwdPDMvjPRgub5hJj9+g0
TwbxGEsB3dJga162hbAEQIL4EVanWdn9txApABQzyFAkaU+RJ0QO+P1p+ou9hWSs
YbXFRjcr19+XCXZ0gpzIkv2Spwu2wg6YizK5P21SPIJvr4kwUG4ILlBOb47AiHgH
yDDJCO+WAvmn4zndzUwJQvL1LmEC5Y/+wnJZ+FJJqaTDRHvCCEPoA1XWQATQ7OZj
NG9evK6iPy+S5TYJ/T2emD/u/81EcH47dJR65wFZlCar2vaL1Kf++b26qcwzPSQf
qMO21ly0gftFm6hnrHarl4xXfzoD22f7CC7sCculanSYHy4dBCEFVpKVRlIDPHUe
tMRDBj1DIJ7Nd1kEZAd2eIdy5nigPyv03m+AbZuTU4u4CNhtuyIAvb5VDlIkMfdd
3glRUDF5TCywoCa2hmYrnJlaR9U94i3HuNttSRgjan+b+q5ICJZV994FWOQjZRni
wl/olLJTej095IPFXE7QNVxkYxFhOsNWBaXHMwNyJpiU2ByPvWvKUEOH1f3Rzb8P
GEev+vKvErFfutjtzT9196Tb0zZCMZrb+BZuXFDsDmmJj795wNdrjFzYna4MRTYb
7K0gse9WWx1S5t3a6Nem96+gO/oXjMEdiCsRT+bCfUvsiIZ0DpAb1DaYYVYajiEt
vyp+BNC+P1ZYtXSY11zE0HZK7YPZ5X1odXHYODiHQWhJTavCeH2W1xFYC8BNb41Y
Xwmwz02avccvNUN/A0x3A2onyljoaAjklSUyidKsrPX8dt2zV8ENXpFrmTuWbf55
VPXYt+HMmKz2fKcBkZkjowdPUwmLbJl567bXEFgtWBbEZH91QYlGUTDm3jcVCZFi
0BbUZXF3wY8TbZkyJzAnH/0bz2WXFbxKoUhLpIAOy4WW0IAppXQRO/xcGBuEiZL2
bNhFsGrE9mwGAcLhg+XwNi8VH3dvfe/GCuEiB+kMhOeEalC++NhaUR2vVjS/Fek+
BQr8TBbJ6Y6b7z5wiAUd6J3oRGm42KnoCQzacRPDUxIG8ZxxYz3pmvPrNqSkziA2
6qwuVwiMG7PLgFrNkyEFvHthWAChpMVSS3FyD04MJhufKkU5yyMEIpQNoB0C7dlp
xyyb6rwQmi7b8AhpnwGr4BNwFHx7sXO7sUHax/0rzYtV5ReSL2GopgvkZ/MxtL1+
+h6/tXK+EEx9izhJgCwjdosYBPtP99cwy+kGWeDdHzLXY2aPfyaBFvwi8QNiVCWJ
0BwvO4fycYHLr5p0XGrVaKNuKNwC5KUsQEB095LbuRT2HxUXs2gsWSZ0bFtL2VMK
8tQ/p5wNp8iL+7rS7lPJuHsoEv0ywqfRxZKyfYJwWup4nwljo3g/fGNU7KoRJX66
7ke+2ydb3j45TdpEs6UMwqHTkoTX+j6ZZIXzhRoxqyrmUqVrnDtYoFSd/q+OkWW0
FRUKGp4hYr6p4Tb/fT0Qo90TyaN6j+V50elU9h4lZEon4VblZR87eygpW/aSQR2V
BfpKCa2+/zcA0qSP1EVviH++4/IQlnzX/mN0zsALm47QK97wp/s2npkCM7LR1Afd
PztKp1A5pfV6ZdQzY1ADJvCRvaFGOSm5Qw7rrtbYGSywAUj1b8H7D85wIsq5O5ci
LqmshltKUrx4sndhQ9hffuXfDbzAqAEDEiAZWHOQk53oRqUiK9Gi7Tz8yHtMX6tg
tU8hKlvb4v9DTkNCX5qVp4a5WdrWNEsdEMDARYGCeX9S/0KoJXxUAekFeits/Ygi
L/QqGd3LsMb39hrlhHrUw5lcKJV1hQO64ISXKuDK/a3OGTjv4PT2kUxgRUUo3jwH
QNl7y8/vDRZkB3CihQXNQNvlnDQilengv0kUIXR3mp1lBV1Uxw0+VtfkrRIPjNTr
Nfs9wVeS/Z6/aMQlgqo1l02CcQN581ZnbB/+rWXAS4z2uFGNdUjV5jyLpIWOcHYM
NyylX3cKcqmIZ+Hx48Gu37KeJeMDweHz9qtSfL8/p48Hk2TIq60fVo1VCz70Zo+c
V9DQyjGhmD/pXq7KyCNxR9vHLDIINl4O2WE4MF/f56u7+f90hUjI7zMGb4F+aszL
84do3ItX6kRG1MFBzlopt7jNqYrYlbRbyj3WUDb+htyAnOm9v89fWgH6nGpbsYN+
eaeTOl9NH/DEHz9sZpHurZHDAcVuzy62RD1pfa36n/7GH8WQnR3cSd3ntg9mLjaF
ki0LMLTCj47e43TNBdpi9HetsdAH20sMsIrWOdSBMpvO/S8jRy2odO6m071tYFyH
PhxJz99iWf0qDH81WBFHAx+Ep7yzuPPDDyQuk8P76N8qF70QuM3s44ynFuFRU6Mo
DKHCwme+GLLeriP27BHHCcuRaz/RT1fSrzu1es8CkxicY9ilrjLjbMOWaQWe65dV
eTktWHvjEsQuDscEAZg9O3diL2w29AoRAwaCSaO0fCHsHax/3kl4PMIWcKdzA/Va
EkNWVhWuE+3qRn5ozc8499VU6TEt2O+kXpy+CdEByZEBUqt27O7lnT7SWMfGvEw9
xuBQRpkqWbVoddLzzl1QPfDull0ViJFti7XLmQluBG776Jgv1HTbxMG/YQW+hoUj
bIusfCLWvStI1nx0HLDJPQdkop0nUEswRW//er2hyUBv16ZRAm9kYTus1OhV5jQf
xjxN6wGY4rb6HTGZHhOTNVmiUyp7ur3g+Dfm7gSslhV5XE4FYqVB+k5mAWg1gRB+
VDPZZTRvsO3RUnhrVtdLSJhjdOT0mWMhSf/LDiEINrWvoJ/8CY97Uz2vVp2o3lHe
TDqA8EOOOnU1rDRHlDPhrVpa+Dtcs5Rg/LjGydR5zVs/H+GkpfxD/hd52UMJLWk2
C2sVt9HsShdzj59P/4mp7gRYkNn5wqlres+V3oq1rFAGH+7h7yptkaK3goq8Ecis
wLfq4/XVSsYbSmDy5dilp9DRk015fJA9CIERWqxLwkaG37hLVe3yWV5QINA6rG89
p1C05WmGVOYuAaeJcVSw8FOzzCX/ppcqWmRU/dS5O+K6uiJ2o6CQ0ajOk/op4pxv
DBgNUzF4w9Dj/zNTkm6VFp2Bp7iTaqaY6hRANoEF0gGGxLn2dyTH5akJaC4e+lGh
SqtBovpgfwKVCP8vo9Ht6QQUbbfLKQ5e585vq78tfS/MGEpJVCkn6IxX8wjy5VNq
og0PwgQZwFotysFwO0fEIcO3SchVhGhqeyUKCK0C128/gEh2BEnZaNga3h4D1APG
onxc1xQfI7AWwS2MElvALXVP+Nr6TeRbc1kJvtFJMTPYQBVDtcGvpZbTypAWO4PS
5aTymWodOuSvVYf2ukOvgRjVOeiXwNybZuG15ZFYqJtu43B7XvO5+ZRsgg5wMrdk
9WS7myjdZDMvGLq3IOgWayPHLTDKevNP8LgTFcAC80LxrTFaVosBKaBTpAtjB68Q
S32li/vdIVA8R+6nk4El5acEUNrzOybGbOubZiyGLxWv4AKwuBp3jucXPHMFfoMP
4BabgvgR8r+prXz7D4O81WS07DqrdV45Rbn3h+UtyC7lOJLUsu0GjRgxq6DvLnlZ
7j9SGVaT+WnUhfUKpWBsHIAHo2nMv8UiDx8sEJVvs9Rg8cGigz2l94W0rerNJ8rl
RVg5CIf1iiyw8Hl7JbXHFCe61QktnqOsX/waC9gVUOS6gLII9u2Mb35CNpI3J78E
Uw0TwzCD1LnmYU0zMtWhNbGlyycGcm5f95MzAF6n9YYRBFzsn2eckviJLrvYoH8j
bT9iBmEMo49ME0QaxXl9zi4cKlsbMNCCPfw+kdnXsGLqOIQT9iNNcGIrOvHMrhUq
0BUcMxtPblEswY8CrhBwQ1HVkFstBmI6uN70SF0IVMdUBE5kmmif2Ldf9ACWFzUH
Ae1MtREZIDADUHGtjHMcKdWj8usfcKYK+AcDHXzK8qNP9voP9SWosv3VvPu7rLEb
MRBXjolM5A0E/iim0sBwGwPbd5QPJLJutbjXacI/a/OiEsfL6//jU9qX76PA2cFc
GMs1eLe0I1MjW77PAla5HZ4u+46Qt/wqSA4YUM5TRP+LkeGXVwZaOD4dPKomDKWt
AahPtaqLJ9mpgDRDeqKTm3mv5Z2EypFf3L2txrhOZKwOXwAbqM7yJsO+8zzLITP8
xdSCr12gFuOm7vf0/a7+gXV+1CuY/J3rm9RgHvaQBZ5ATNsOA0kT+wEYtCBKD29L
uMF8ktSWS3MofqCe2978gIocipq9WcmEY5djlKfRNI7Dq47RFg1dRII065RZozlk
xMNjMfYA57NQ0Hj2iTxujQWDcyZc8fX20lc1LwcPsFJzps3CnbKeptggyQflj79r
f2gFZgADJfrA1B5IYf/l0e/4gRsirpe55PbZDx2wmd+igM4BlCSXPBAS+PyJ5Uk0
FwicjAeHzwPEyNO5ZF5CCgCarj+mEEgn9Ru/Xe+ndUEeg2ql17jBxz7Smy5OpABV
Ns/5pSdfB3gvHUCjUnNHhKEJnxys5yJMTI8kKFBGKHB3EKaGMQM7B5G4QVRrWHQ0
KgHIuRSBxdKENhAfR7ISDJVOV+RtYTwC797GVEfVG7Tn+loaFsPNj7c8Bi6cHeuB
QHUFfiKfVsWgi3D/FyYkq8sKaTNgFg+mDeUE95z6xD2ST/bm1G6yndhbWsMX1US4
9+oTPvUbXDlhzTMFGHazEe1DLTtIW/9FPJVxWpW58CFjsEh/XGJSxag4W5Wcu5Co
Zk6YSOxEoMzIgmARMlLvxpPUTVGonVs5BIRGauLHFB1qBSbUhmweL8pplCS2tku3
Py3uGAEaxMu5kOsZdoU1NbHhW4bPsKDqopjdKKEfUDAoeSMKfX685Ee3fCUcwbrD
DPEZ+PzoDD6DsguVoDgUlCLl5Bwx8tobn2fuhv+V9XrCQCB+tmYxWyITqBpItdVP
bRwhpnIBkx3snOdnth5kqVjc/+5GDonxUu28NT6j4vEr237hdOxBXs8+btDMvvBP
7j7xh2GdqhZphUn1RhBprnCGzimtptdvCjV+bIxuLj4+IsyH/EBnAnyvmJD2dIZl
8fY5EztrJSs+EKC7OewReEBN582BDGJBJ80xygd4xUTCBYVxdpVnkW4ddIXW23Pk
rypof18hDJuwLBGYxuNb3gKZ4O74DS5KEFZiscJRSweLqKCVJm0qLljLtpGHli6R
6WGHob244bp1+lqGQ23AEhfBxJOfgN+UszsAb5PE39rxi8HrOuTC40yWTEPVlVPs
VkjtX2mrruKsM2r5PYzh6fbLp6qkaf7CKRN7O9XJNTzB/jfJmpHwmiwwvBERoP03
s6DaTCPJerDiGXDVGLgDH7xn9h3cRvOknuwpwkqnm+GsxifyoinOoUJriVAx2ESs
50VtZBrXFZV23z+wd98bUD4t5XgZvlgFuHfu39mxJJfHpvJC7qu8n4UhI6afAbjX
RzQe2AEPHYSGyh8QWrUja2rSb0YMM6ifjSg9Nx/q2gqVf+n7B5UzMpXyADrHJET/
LOrJ7an5CWNmJC+LMt9abNOwusaQqWqTixgVk9cyCo59zdR3uHXBs8sNKWQvy7hW
yvFtqyP2+YAuBzRUcmj3dZ9VCXOp53GbafjSvkgAPrU58mpFJYYxZbTTice10k7S
4Q6vBzeuEc0msYMbqwnjDuk4it76TWWjToMOqN4vcsfeb2EUE4UoWJijYRH4vMHt
P6IvbIF2087s/Z9DRh265Pb7McGkcwQCXve4/Z2VsN5/Gtp+82Y+PH8CWJZteSIT
lH7F1tWGffBWtMGK40MBwcArTbjDoGO1K9FV9IOSYcciqs9vTqdMtzdY5Sh/PK9Y
z6Ik1OIdSt5Ba1jfSSMpNfVgRcG018j99le38Iy1cxSpkln8mrC4UzDEmZkrJa7M
CTHjRpoidC2BgOftrfLwWUytyLV3ng3B7Mn2tQyi7+3EN8sMfX6riFm6fdRG4XQr
IYmspTvep489fFNBHaNmZLzzSIH8QAEY6lXkPtJup4ulqJ0W5yxsSEtAelwZHc4Q
e1huq+jR3MFKFu7eEqa8pbaLZomNrzxOTUh7/wJd3VT8Nq2nkbiT3uCSdKaKnofa
8ARn/JdE6GfXm5d7gw+69NEeG10l2QYxW/XF0Dty16tObmEzJ1AUR0hyJIGJb1uO
4I8P2VmmCsQxS4TNCZoOcKKbrmboAs7yTfWtP4M0vSeRsbqG1ULu0T1vOusiHrhE
AVHd2vsVATu19DMXqTkSe+xTHJiULN7R5kkux8jOF187aFsEs0uUihL1qtKaueLH
wTATjCtAubs1pcbG7jHLx+EzhoG8WF+X6V0Ol9VCLsDcm8YC/yMSuQ4FVHkyKhOT
mmhuyba68Oy7T/d7xmsheFbU1g4PCyrqh3WlHOrtLb5yhZmkkquV/XcB0fXI877T
H+UMSAYZklfNkXG1joJuWFfu4+jFs5T9LbAPMothwK6HoxBpQgQw5TGVOzQbeIb3
/LvxrQF/Zrc07jY1BWSMi5lK/rs8sGeusxrvgVVYqkSi/1uR9Bec+ki7BIbVi991
wDbKxlb8SvN96skZWEDbUXVnsGeCcpIMJdbpQL54c2pfqJucnk4ugbDMorPnTDx7
QmTOYsSXK9PVJuco1Zr133hyapC8rcXwfohopI9tKit/o9M8Zsu1HnBQ5M7EKTuc
k7L+VDgd5Nb31kzNF2OHDbVlA4Hf2dKDH+nDUoLkop4irKRpf+8L97xou+DqLm7N
Tv6vaqrJrL1Pf8TnJ+o9qPrBlHElC9ohDocA/2mg/xxZBZjYjEYRe6JGc/C0nsfv
umK3PLZjO7vtr3IENwxdF1woxqLxiaZVnXDrljbFqZFR3EiniyiWupEoDZlMbnOt
fXPTEfcStJiOvGQlto9jPmN3nECHQKuOslPC6nJRTVwAT1l+H6OG7Q+KYKe9i8M+
hEPRZRaIjq08/DzfuVMLAi9ymW58/1JKK7sqf7EJwueJg/pDgL3yEBvC4rKDvR16
EZ9G3ewR93mevLKAehaovjzzkS0lbQLZvTMbCwv157JAcjA/lL2cBsv9H4FKpHiN
RwiEjeGt8RFDXIx87qHC0LbFe9+zY2PJkn/doIHyAiTo4xK9fPqic5kgqUm4/SOX
bazGsgRPZN/TDd/9mR75097z4dug36zfjkbiaAfHgDTGhheRRMe5fYe7BmiIV93w
71t+VhnnM6w8LWMCHm3Zcb5XDBPhvvZ0ZAgKvonVaIfDU5hbnvB8L7KqShSY1pv8
NX49qDBFvYYbEsAPgFQg4D/9FQbcpBoBnHczFclmBgu+O94g8ydml2lAT1VfBj9t
Q4nrSi45SCghL/+kjD4tOfIjHN1pXTTaFnSLKEOBrMv6LIY/GtQOD8z8r61/2R9g
QvLhd7gD6ybcES5Qn6qTo3hrmG+gvm4CGWE3b51PH5qpdomquoJtxmQM3ATIx2Li
FXbkEhl+iod//nZBYkeXdZzgHyPUsfFTvvPjdLKWQVWjlyYC+do6MtShNPHVRBtj
2s+2I1Fk1iYix6tknbCoxZnV5zeHJaIXqM2hjMIS4kVSiuOVRCR4tpOuzCNhtoo+
BqWBbNDynSsE1VaV8sFosUsLF9cDQMd9n+vixSLj0SNCO4EyF3Ko5CrsthMwSj38
vhTKjL7WB1ZP8jiA0PA+mTE2AQWGxsNiwNoA+F4fWdicWSjp+68u+g+3l8HPnnMu
PsKXQrfrLH8yjuIfSfSaabrM89cvb6mMy7xiXBo83PJCCSNAViHhk4Q+kOaTgIBB
nWui93y0Uln/ggWvI+/2pr3GNtGLEjgNrfTLhSmw0eaXi0/DiJXynuDXJYSK2JR6
YNS7ylqbHL4ARYVcKcwrjOFWL+FieiKly/qsPATorSefYt9XTbEPj09FiWYBK51V
L2nhfD4iBYQiPoBb5saQi/duVGP65A5XYwb9CVcpkVyiiv2eA/Pt4T/GQE1EJBmq
y4Tkeo1jksG0rMsus4qIuJqtSigFsZZKpP6oh1upU0NbMod74FCmp3as6g60ZDUD
5vmOZKRhE33S662TpGz7NQUbT0PKbMDNUJMv9UCyhCVwgfbjuh82zLDdDZfEugPC
G6rr3aUEuFw5ca/nAHqh4B57QXvduxQO9BOFWBw/AD1aoRr4UHqBm3yR7Zio2ETX
JV4MaeA9xdEbQR0a3EUOdLJPsZxSFABRzdzu7i/EfNuKrSb2oud/lAHhZYMIZS6I
JMmo9eREiadvb9Sx9q8Txq+YwtqoJN/MMjNTMpknpDO4Vcyt2yKX9MACpH1agi6t
q4Q6UYTjNFpM4oy4B07wAs41cfvztTrJYQfRn1GCVbJZl4lGT5I5fIVcH5lejD6Q
wRrrvYRT0O+t+AAnerJG6U0qlLGxOj4KuNP60rd9pXjl3w/KhXY1YoSicxHCh9fe
aKNM+2fC+jpJLNPpVrP8qMX/FXEqn+FgYHPK3NQRLYJZgQRbHNiPTR61TtWfs50n
4jy/Rdpj91J+3s3sLVkeAidF4KLbB0KJm1GxdNyf9MFk/yz/AKJhh2EDPIIeYTvu
i+1QlB5voUTGAi3rFWxhaImrNVK7ipU9fr2+wauG2FVp7xl7jSdMwbalbkI+w1WX
SiBq+nwnKaUKrUs7lNyIIESOzGnXia+fDAnyY+nlISO2pCiv/1KUdRkmQrL2jSht
lwC6NUTvo5bl2vIPH9TwSZN6mtaU6fmYeP6tvjJs3B2oqBUT7/jOhlilerMTcZIJ
IyJkL5LgQ7j0DRJtClj8CteQ66s4RgNxj7gBLVTsCHA=
`protect END_PROTECTED
