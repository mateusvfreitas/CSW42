`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Q783K0GSiN476ZPh6sijrt00pqH97XxyR3UupBgq5Q3PppiCoqvf4H9n8ebt4dDj
8gU+sfsHT3/Ju7OW55pHnRvLzyddZ09LaBdyafzzT4cFi/tJt5HOI/Y8SoocK6BG
D/n+lecREnDePpPhmBKmsi4lo1ssQ7TWjP44B54t3egyhwXgIVeDXi1839muwGy2
HSBGCTi84OJWW8sF9TfWlI/cxR0s0oP4aeYDd/8kKUhgvBLXcPhfAg89CL/m7Gkv
4wVamG9i9MnB3OkMulVdLrKV2ZDC94uqG09k4qHI0iaxHxbrrq2+cmt7Vh5uMRsJ
9gEzn+LU+o0DU8uHJ1IcLVbLk/C/c85vR4lY77hpyNGs1iY/j7WbIgOaexSE2cDm
xJZK53L5GyWpVREMgKxGR6dJqaA8xVSDtZ87GsbWIv4E0tTX5I/QIuLV6fZzOm2i
twyh2dHNi8ARCajOxu6Y/3QBF2lPTVSwg4tN5naX190Wx/9JoZE/TwUWfty89UBd
jgeSgcQTxwtrbSYBHcSNsvPnuQTleZ73NbW1ImREZojOf8X7AxGZb3I4/3mw1oqt
vvIpnmlyGpo/LQEB3QhEjTvnVMHqn2Nr83KdPm7UiqxKOeBoznYg8cCLALbTlYCM
Pjcfo/2FRL0Ge5CBSCxTws4lJ7nNHz6JqQHVyUW2sRfcKP/hlt8MlIpBfR8Mj4G+
HYM5DxKZmCzlogUVLAVR9qbBcBdMG1ZmbEwtMfSzWhnfm0y9ytLlzsU+/CFLCng4
7kyuRk161tQjkMcHraJC2jvQC0DRW1yE8SJ0sRRPCEoTDRkH1zNJBt6pSRF1x2A5
9iACZrc1giSGvEm6xyF7Padj3+FGZTWvx1quenAqbdGiLU8lPPvs7O8uFZYMquSl
kTDoAQZ6ISOHK/59lC/T73d3Q5DRyGknmMcqfIV4MH3xp68A+lXjwLiCwHq6DnmP
8rQy6topbSeF7fUtibJvSdFXngpesp78lmDoATXtI0fsv6BQ5W1QrULU8je/TAuK
23qDYck8odN/xRKcSqIWnAHY6//DzF2xKhnfJYvvNZTmRNMYoUwwbNRo7gqeWMmg
bhyDn6RMfzV3g6nWetLacoHlpyYeT+pzay50Z1Nr4PNtsUYvF88JCNsqYzYoxJDY
N0XMXn6tZqB+v26O64K83w7nFItZDWBVGhnVuGe7bQ9rTLurt3XMWyw+NjD3gEnL
b32wYTsvkB7pkjks75IDVmHWmQayW3MbcUjW4D1nSigzixBINUDjknpTcfFQuUJr
+YBiUapjOj5mpfIyFy0nV7kULM2qV5KBfESF9nyOoY8iqgnYVO7x6R7Z/Vaqnpgh
8mKC3w8HiS72zqx/Md6F7+MbguDQv795L9+qoyJZehZt5CM1+UXshN1mu7Lya0RO
CgpH1b7tyEVV4aym7HBdFfyXuVDK27jU8Aadj6tk90Gews6YSQfaObAvtPHvtBiC
qUxa1fhZMNMc3ZmNyDvgExCugkrBuNYU6T2/vxffAw0UYMtjunCGgWbkLyuFORHF
gplFCj9GI2/7fLSDV2bsxpBgvnAmYifnuYhH0Ta4NcDITdeXPkoCh5CPH8sKjDVJ
I+HaM1CqKwmTvqiZ9KS6AG02hvQUwisXcTFsjw6m77CuQlFzdWAVqxddba9bCpX4
PjcTA4ZGaGnKieUfnUCxdCecT8K35ff6o2M7lBs8t+vL/8FSr9AuynF2m4ZOnVa7
nAdO25jJcID7atauRoL8BIjHASw+bOZcbRMnGprNpXh7CyZvM51Fi5ZOYLWYDJwl
euMkoNJw9XcWjTc+ENyCubiv8obi35liJWwnEhdWdFXw+d7apQ1zvu/MaRV6cLKC
WNtc0Gol+Yz460nmMtEX8/cpNa05DsMVuJ2iOwa67zB1ZTDU3kRh0kiMA41wHz7X
4OcTU+F1GCEsbZu9MeY9t7U2r9cufs/LnoVwma+Y5RqXMNZDCT4pnd8g8BNP4emJ
6Uaa7opUUSt+O83SvKITousE/1ZnF50M5P2pgDMJ+7Hm2CnZt97UydVOuMEr8UuY
loGMhMH6/PZSR8cMkVhK27uw5OXQrXOl+LA6gJs756DWyxv4HlgJHr7Vb5+/YQbM
+y+QWmPZF6MLxLOcxxl9vQxXE0vLCJZOvR7xR7B3NOFW4Tm5AdG3YYpyKpsD5dbm
OnXmLjEDbA07IneKNICV5rKtxZZOWgeQXjVojld4C8RkYBTS8/SvSBHVwlPqwp5O
bWemxtioyfVfXHvf8aIDobmRatlRRP2cCjzv31Z/Q+KDIKz7sCb8ciao/UaJogKo
KVs6AsqDW5VgGYqQqU0PA1Z836vTzbWmxJK3gHDytDqMcuILupkMk8AgjwfMDW8P
BvhRuoh6LlXpFXDz+Tk15l3mUXlKEXxcJbbt1By+AbxHcWwyB50MHu1v001FiGIv
BIvEDkwUtFN/LrdxggExX20UAGgDPaLEZPW7YTQ2pfXo4H5xPTAaSCCkQjfy1wmg
1o0lqQeEB6NgOYUwFghPTXzJGRhyYMLY7PF6xWJxTzC0t1D9iA6HLEUrq7L4891d
zlOLL1mCl8XN6uyLHGqU3xw4rVGPswE/i1hTO1fbwQD3qOabOjwPC7ymNJ+Veoct
zE6TU/ggTEHT9iDDtcm+isiaJNuyZoZIS2OwfHsQOyMGb/oBPN10H0ppTzXJ0HdG
kXbASLVBd1YshMydopObGWjyuT34uD0tAbBAbrSdIH8wdZvB3IkRDCeba3uzbVFU
2EyBZZHYEEgtf1k+wRCzMvtFMEYWnyrDkdwLVY9WKNi9WTdB+hhqo+Huz02/dmCb
8MrmSVTk4LCDE73kEkFxK7isy3tMKUQTPdzjk8+zAy95i7xzkMcwL5C3tC0JBdra
I2MKB1drFPvwxDxEHinDik21U/IrOe0fkHHQ1G3X+EdCgUyMq6qaDSmpk0y2EFyu
74e46C2pjYXTRVyYF9ZMyFgPGl7J1iEF9ljRB6ofFMtuL6glg2O4xce+Aw6DERS5
lav84YPnOKdRg+ks82juOu54rnyh4GUViXACH9flOZiC1e7KDd1NIaDrjbK9qb8B
cg7vP0LhWo/OUAJdbVHcSKHpKNao0OnH9VDPxPtchs85L6v0PDMwIZOad4k0mK2W
t0D9ck02Bx9Kxwq+LCguLLDX0pE7LyL/YcXAz/PwXwyDkKrILp8dtbbtfAkqQsOA
HdswoM8aAoPN7Yx5pgDwMaDwhd3TmPGlpM3+/cvfDOG5Y5D5fLY5VNqpd8R9HXlY
GU0cOVceOXdzFsfUo5pL7QIiuhZmBBe9hWiApsTs5oCKTXOf3p1ZTjiI1XMN/Xvt
XpqPPnxNsBYSyP/Tgy+SahANpr2vG0b4PNhQQVHDw6IDpey7GdvWGSR13bHToYrJ
hBm61zXueERmeLys2V5VY1J9vkJ1V5R3axXyEDpFJxthv6TeB8tJdHGi/neZCQQ5
neu2Fk9a21TvngdBdA+UC1u9a7DfaaBuLJezAVOYvqbB5gHmF28o2F+M/bNlC8Zx
sPgfJN3Rlv6TJAaIZyyA58/oWs6MAFlrliwTRUMoybxCQG1tDn/mIh+RHLmdLtnt
EmigJPLbo4kt9PJ9Gd6kgA0qD7VwfNWvwcKxoC5u1jXa9jtHinUoCKwzhbiSqrLR
t6pPFHFqUVENdCnlhDsmJ9ruG7djvcSEa2a/vb1wnS2ew3PSJ8apZLCAYzj+VwIl
ADBF+eSnzXZUn2+r1HS49QMN6iMtr39VSZ0KNAYc80sxx82l5EA9IWlt7z4V8kGH
oaLHTKRFmslNMB3nVTL9I9Rq6Z9eQZs30d/vYyY2Pirhxc1nmsnY3g8TgD5kSm3Z
T30PdEDWIfUjl7kttgwNsvwHZVaxNNNxaD2rfuGA9AEW1ACCi8KnK+PSRxAfnaGq
1uJF6euu9s5dlt37vLBZhqvkjfqnJZH46WPjmHNOl5+8MdadWjq4vCgOKqigUllB
UzYJvBG6c6Smu7+CJKrrQ9TVZEzYY0R8m+XrbZQWNVZDFcPr5dl7NdBM4LELClZH
QlsyvrT85VXXdPthqGSMzrtSO2RAC745ih3nYTzqJ7kkXAPB3golJsE1drO83wut
tPO0ghp+2EfD5+4oqAMRdNJcjIFT4l9mzpqwdiseGhtlo5WNb1+HRjcKYOxHJ+r0
cjXMJeuxQdihUGDRWbOivQz0tIFqleOMKvzXwssS7p2sgDxGC8Pc5EwSZBFHz1w2
rHTc8KXar85YhV5GHYuVRbkfxACZS4ZKsGlAWL5BfaZZyxYyXMN9//NhF8K/w/yo
UcWrJouZZByzfYys+k73zyEURy8yVsLqT4k2kP1tddglBY41aka47bqZzUuXK8iT
eZY5M3HfepxfjAAWHqZAswu16SqtgLHKpnXmyQqsq8wdIJNtOfFlmucQ0kaeCMCi
XF7JyGJMUzwj48bPOc5sDvwIxwqVRg/jFEALy6UC8caYdesIx5/1znCIpww6cWMl
rzgEd59/m5yG1lO513aYfMC/6IfIG+rDCYhN/6V/TB/1LTM4fciTDBEaDWkEmH68
tjMIp0bt2DJSs/jUJKENKqJUxp0V0LX+yqVHQei7R6MD8Y6w+VW9wFNYYN5F41nL
PBkfBzO2M6WhvhHh2q34SajTDKOK0bGby0haS0YmS4Y+QIK94TCLMcVI46q0WZgU
1Vtb5retRNl/8VUFifXg1XnK4hJx9EGORD0Wp6ja3Y8QrMT4EBQf1c4a9sHFIDpU
jxwN6cKxs2RMXI5kz8GRrmfg9VLS5iFrVa7MFCbvDJF9KQPq8nJT3UBPDkEBhDPB
X8ejULrHuzRbiV4K0XrGd+gWRNCmtCEeW45GAvwyNQb0VYpcAKFLMh8UmStU8MAr
ji+wtTjuPa1/SXqKBcg+Y9kkpg/a1/zpczT/LBpD2ubZVjCtoerxezQJ74Q2VR6I
c3ct4whxjjds/ZcwT0VgQGb5EBHhzrvkeWEtcaqihMgYYnUIgzP4pj25rD4jsb+1
635Xqtlha1WO8k8iRz1ZaxQeGKMW3ebVkEaT+vpKgoLho6DET1VYEA70p5UlAXJo
oXvl8O0iP2GX5DDH+b6WFiTYDidPKOZ2wobTJSRoZ5DjVZH5lA+jLdj8N1vOVkz/
tdvt91BBs7oQEVEUZcw+KHpytvXzZJYD8P9wIc56YTMac0T31CZTKoP2mnV8rYXj
3VuGn8kMhPLYeMjZHccvNQrhhbAUaFiCtPRVpH0gQARvvu7gZBUaB5Fos6ZDJCW/
dkftz6nAmwEdNRS5DPPhMuXT+76VNKPS60wTKxpQI2sPfS5HwvmIhV4ohi8QYbn4
1n9tucrz6ubZSRT9JYTV6ZAJr/fgX/uC8vk1VXK4d+yvM2BwOX6h6ENH9OMQ7TWH
cbJvd8bG3i6PkYWlUrK2OI4AncxR2RElZyalH2lueY2CJ5R1cczq+rsRjeHQl8Ns
2bSOZQdF/3rT3g5H1dfKrsg4TzVFEw4dIChUxEzi1r7XRKjNdYTQGM7L4Qaesa5m
fxrbe6TMu7zM/mnWx0zGTHsbyNJtkscoA1v3P5j2A907ftZaa5jdf87gb4PGo035
us0rkETEUCnWyGGgJwq9RozWTxh5N0334LXg+zLMTS9SlNwdIG4GrXb98vrMeeHL
pv5deS5fm5bEK8ZhAlMqLA2M3gRltmCzviUF+UtvE9a/0g7dB/BLIwYXnckO8zsC
cZsvYBktQtzyJ/LVd3wwnfehGQFLozyYM5FwDx7ssMHv3+4K3p08b69ehoOGVjW/
MCSzqXjC99YE70jf/mSLEabDAEzPY5DU4M/L0EK6+lGPFDQkx08hr9x7t754HYIL
lptdF7AYRWwnbOZiQBTt9g5AQFV/EdkFe5qaNjhjIQpe1gxHwAaBlUSNdPaUXCeD
fhojI/Hzvglmgh27xiXAcUwXG7fNTM9DAWzXKpgm4ytIOCM8I/Dqpwlh1iibnCj/
57dKiqz2q3+ULvxvkpVhnlfJYIStgf2ZbQmlIMLDrXQ4AzbpfYv9YHkR4daamMab
6xdzppC3aUjwtLw2gxw+s1B8x+9BzJiYmazADN8qShQ=
`protect END_PROTECTED
