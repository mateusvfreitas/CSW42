`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
wwMC9k/HxV2NnQPA79mhDS2U3rrZf78bVMNs7GYg/d+VbkUS2DiaIBuv6QhJQQwK
0+GRgtg5g4j4cU6y32WwYV/FlQi6LYNvMoEBvX/mifdI+Y3SiJJhe7Gkuuhgc0yP
O5eUUmTpQg9ii75mzWHfXacLCVNYrCbnDM3RWR6fqvRwv1zLYjyXWshLxRdtgSWE
074AcS5P7Rf0L4VzigpXQ+GT+/zQfdTbbLcsQFO59jeUGZnqgROtvFnJEg9xLKRt
ldynWdjSeXBju7GbRf5UfZMUWAqAlbmiju3cmpDemKMZJi61QmPzHA4Lgn3ii9wk
7Gzj2c2Owlzv86u0EhhJDBITc7NxDBjkJRdrCc0vhOR+GJBd9idMW6VhtWSnYPvj
iBPeyoESdWPY/1tQsOvSC3Vh22TiZwVNSaQOkkI9NPG8ffxm3g4CIg+kK5gGfUGj
J1BPpNtMQQrVKUC01N7Y22zXwZodImIP+OcICrFSQeQUPm3uEJDMnYvzCLWCfZaX
axh0NVEph8qMdFBcj4cgfGZPotOHV6ESUVI1fkSg/38EKt+WagvHXgvgZCmgFr7+
9ErMSYzeyUuPj8cLe8g2HinU74uAq4cgdCcrsKDrvGak5RXflZuS7SzmZZ+7URgM
LdbTIdVW239xGm19f+YAcb9gHO/7naPz6y87rg3ixzm3aPNXI63AJwuMj8NeQJOc
rvv4Ma4Sq833le15T0QHe3BecM0cslTsN06npfXZ7enT/Gc/EcFQ1ar9EzLI+YN/
fCEO1dzJVmPUPPO60Qcbz09X0SMEIFIQLCw9IOohe5dI+Par8kJL752/kv1ZkUYj
bCS3/UQnHxZIUNkiIoM8OHDBkRRXO64R4a2Sk4rnVsPw7fdiM9+VTHt5/F5AFn+K
Jbbu7Yh6g/N3iddx8PRWdhZ7CJQtkXybXQyKCAAwa1V6fmQkpscnnY2basuQfA4j
XTpOUrM90xNSF58D4YamquZMQGiexSOd1R0JgPcCOzPgU4zJfYnaIqs65sPcRu8l
UfO5tZr4Rinh26DuGwJJNeqep0BkmKbxRcGNkGdE/McTkseFDDeDsLHYthdF6RaR
oNCHP1RO/TU7mMehdTcj19Qq9RFFG0AYKkB71RWZtcYK/54SATvGFURThy29brl0
VToXomIPnFY5iBxGkK4kPo5zZGbq2fFcpeyq+P9JVqKLfnp7CYsAcnlkvo1Qz85n
EwP3eeDoW+Ob2lojyRvmhI7ugzk51Ep2YUAlzxn7lASES1BKm6duECZBl5L+5cJl
FeUYePnvj6u+bNJqQ1qBgckGhuIvKBooQGTByEMK4mc225nHaQh5tFEWg1L0JWcj
sL0AFpn/OjOB+TUCj0IUPuBYc0T5L9fcPnN7inV+LZ51+9HY+IFeFq+QW6mPTtO2
zZStyXWjw8XNrUO0QNBVRNXAy45C2LZNn5+QukkXiOJ2nnscajIUzFcN0jyhg1UQ
35+XVO429zb3kVG8RVTf79oaQ7TR4d1LAqpL6rb6eKHC05eQalAsIsGhJuGjKi6h
YRel4v7N57BK4VPQpFLbynHHOE2uXnG97pcS06It0z/VHY7qHKmseGn+X99AiwkW
102S2ZcaD9RofIlqEIt3x2IPi9FNdViL3vuwYNj8bMEhsksE+sch5tJBnrCZob3f
P2sRysMhNIpGIku8DgVZpWX7z4q/IKDFVCgX3RyKgWgTSTBF3MrWbE7AnpZYMScw
a7/s6EN5sKgY/vBZBmtDxRJlqnHYjqipOVUgmJUimQ9AtwAVOAFjRCu3Pxvz+e6N
fle0K2wKvkAwSm2KMChg8g9eBj2gvU3s4xMbVOI49oIahnT8uJMf8KQBKUQKh+as
CQkiU6+7Rfufp2qpNfnH4oQVaUoV8o0f1iY8yu3TEJjSAyX16KYFSSsDnNlIMyHp
juDkvS+roYFpDHfGmoop4ytaKMuCLYrk1oCrwjrLyb/vNObfG0px4Wjl7sgHqomA
IEFIiY3OT/mnhs5kwCVZNfjNZmiJNL8QEtvVsLjtDW3nXO2aYPyciQNNKwMnijCN
Woe8sIJ2E4gZnEk4U02YoSqbZoPHORFR1i2uDvCAAk8pMoD6qCkmqsF9GJ7vKulj
NRDYpNGI7GJz9rGWUMH+3u63DGlTFtbzCzosF86Cbq9CMCa3d5nGVX/6jSCdrM7H
h2COpfwpld6eksRUZdIY89loHhaCbJbHwMjzE5opxcV/8mvLtWpEAEE2FAp5zDv7
LIX4gK3UL3GFTaVUe1iN0bXzLwTvajNsqFg2+KMZBr1AOBmKBZUGIT50acPJfLP8
kiWDbV7bgMpe6QQjDQpcyvC6/hAdPDEXqrX81HTMGahwxxUnC+gv8S0IcUR1ZzO2
2nt/PZFY5/wDh50e3fbJVH2durz9YolDKxG0CRjbnusEEbr+O7iFNMOFFrFRgTIH
KwkdtNRPGng9jHBqXItaBNMXY2h1M/iVi5iqHe07DVinkrVkxPCuFruXIYo5DurO
4geKk8eNQ3Z7sWOxabmTbyI/F7KDL4pjtqq5i4zonW8xYrtQkSXsyHOjXfguC+Oi
9hgtkk2Z+ZuLdKcNNYULvTipHRPS8ImR30NS/4K5qJ9uzRq0m8ydpFSC4zSRUml+
G2pg0b+6SfkstL++k6F4S5Hkmoye4bFHoSVZ/Xlyu1ocX/QXeuGBfnbR90/jyAWO
JwAQEmvRVNINDvWgY2EObUbamHPLBJOYzbUUIHmaKubGH27z99w3MyjrFGSIC1w+
NbVTgJ3ope046Lgru6rIeA/PzEHgLpkV7cJRsalSFtg79KK+xR0VRoLj2YCOd22d
k8M0G/OGpHrwT3NDP8d8BWPMhzoGI69gr5cJQQB8a3sj7KTdhpHugWLgJl0P5Eka
DU6xbewUORlRkuf7iH0a58ppwi5VV/Qr7+6Eo+M1VpmENd7PGcISYSzISzj+8AgI
gzpXJblto/amhUIisH8AnhwDmQOwHHGBNGSGxQHDbb5f1TDLH0e5tw4gCs31Smtr
ah2I1bjxeipD/KbXEg1CCwxHI2USsF+wX9/uHnkJMcs6smui/4zmBihz0G9P2hdH
f7hX5ieS72CJ2x9B1oSsKEqjOpU1GZ3CrOy++ey+Wnhc8K4J5YK+uciI5TUogKDo
qs7REICUjuCIKhE0KcC2wBqYw1t64Yib+OF/pu3qz6CtGRwfn6CcwyyAyR1qf5Ls
/deo12O8bfNMdZCBWWx4oBWglBWgSD5w7lf4/BvDI0GmWVp3LYzWFXdOPAKfqO9A
+5Emydd1Hux9Ww3yejKF+gltHS5POuJW+xrDlY5tBjdw0pLz7HC9Vgs6vayVypyl
BpEP1+R2wf+QHlNkPUH+5SvYurbdN4sqBOND8SenpCzxUOeINstfv3xmw8Rctlou
rYixZGVaADQy7WcdqzK7CohF96ej+rlUm+Vev/WLjnpvVlsD6ac9PGALnbTyl7Q8
Boh9XKpojBw4Nfn8Po9kCNcykJxIKOaoopvLAgsBvFyUeSqFYj0jrAu/SW+R+KGd
S8WGksWS+VyiCsdGwIvbI6avGiRpU3qDIQk4pQXjGxshC3r1rrjIH0co+lAxdkZB
4ZX97FY+lnVY9FUfdIzcqacFkbtn7Q2HIypFS5c9d1jI47nOwSl/9v1v0xV2gCh2
5mJb38QtGL6ODDB4mQHCGDSN+n9S4wPUKawuo9ai30x7jaJtM31nkK1IvkywY6J6
sPNrLolzCk55eNScg3R4GR6oBd4D2lxX7Ttep3iaR9mtcrzmRWeB9+0Tk4FkcpVF
ueHTyNOai3x5/Ap1bRpTVaRqkHNq5Kry0tLkIrO5a8zSMw0QkAiblgbqcjWYXj1w
8rUg8L3gfA5740LpWCRLuKc36WZHNh4LvGvSr8jvOcLtBAo6F/r+g4Lvx32nxwtW
IPgmLu0Py5/IWUaLN6fgdSlJmx7Lbq35qVSWZeQB6OSeN5tpw2c8nN3E/TB4skpU
d6vx8nnnoumOjv50nSEXKjYwkKqWnpCISQU93hjyPKc6HVouGDDMNbV5hgRQKJIY
elpvrrPZN7WcE9uJDPm4SrnpJ9g/iLiz6+DNVxMO9JkUjsaCw9VpEai3Asjk4iPq
mXvc2VfIDbWE6xyd9ykUecl/2a8naHkquo6PYRsbo9uqbAonCcIZS9Nef81bx5bz
m1ymPCuKes1ZHgPFgDao+/xdPMkeZRbRLAXlWmVHh3D6P33XwUU3jYP4tDXFUSQ0
gOKxxLf6tT5PZwF4j/IfZbskHmhAuf4Q+4Euw6AkvQXqpbkQ0VO9U66YVF1X/wOm
CKt95dMT0tMfoxbh9FWcihTIkS4nhaUKrvfDHvANkFSVdSy+x5LJ+a1AMzxb7/58
B7jrveXupPX52U4oNuJ33W05ecIWEP+ueTpjiNxS9/hLrRaGW6iGepi8kba2Ldcg
d2Qf3ZRIByoBoJpu2hx3VCC4nFCNqfLYOydbTKWv5JH1ClR6aYOFzh+VI8LcUAsQ
J92B5SKnjRchrfW0Ppk+O2E51FKucuVN4Qy1DUDG5uq526pxrZ6zjx0rKuIfr00v
m9dXxSLJGLGWGe+XNOJo2h7lZKWCGs69JID+Dcs2HqzbBO4EVWFG56ZVip1Byq7/
EEqIBq8d+NrWWDJVHd57M/GGAoOEiUFFw+uGWn0lXSlkaP6Za0ZRm8iFzp7m6TWM
bCAUzN2M+mJiQMLvm+UeYcGMQAAs9+gKBxgHzLLvDHTWu5lKbjqVOPr5y6xq5ixO
/3eKWb5WI1/EDuGcaneJxwVQ/acZVHCttAEj6W5HeCRBpRBx+EUctbrp/kHYMb6e
QyQXu0IbzDU1FclK2w6cZ5QEqMhr1Yvw59H5P0JBtrd1QUhKxRnwCJaxwU2basE7
pSzEkGs+Lvt724mkDe+ZwDiFD+4aCbRQDDCWlC4BnePkdXIGWqlF0dFM2CjTUNbu
U/0yNIEpS4wMYAOpn4uI5KEDNp2103y6Nau+pgNx9bsb9t9Geeps+B80mM3dVTk5
0hmAKpscRiixfXQXc4gG5JzwFKLBzQFo7nkmD0v5FWSKb3Zfephm2+4ZEK5kaAPV
P7HRg5v5iM15tsbJ6IbCnZhZqKvDV6kuzh0oYEybr567qqcVB8aVEmUJsKwDQvtv
QkxQtBee/djO35J0IdteJ+pWQxiH4ftKm9qLaa1ITLaBLmxFlLa1vMEx7SN/xyh6
qjGB2CIKEqri7lFsv+lPoiYx4tCISdgU2eja3nbqSGu2gTzhGk7czpjpHri3FCoV
MsYGQPT/icdamIAoinaDfnySgUcSaSwXrE+IgIVU+mT8u6QLUvtF7TgstpnPF3xL
mewdwS8iNxR1wnyLsYWz9qN6FAqUhogwAa6DM1m5rtWG5J4nvvBGusNZA8w17G6g
UdONETUnxxveGduvjlOgZmrr/Ww6tKQ4mQw7InXvUSgM85GwMrdtHBxmVn2EK2so
PWhMstbzap+IdHLWOc+Dxy46BLfhAk50PcllB1YlNfvyQDXf1Bw8Erb0oG7jdcmL
/Rr0wqty+1uOu2sduwbVlBHPBV0INAIBPXvOcjqUMe5msvEPBpv3j6SiY3pYSFMV
ROlIILMsq6I8Ot2s82eaLQ4qcrM2CMvFBq8Ho1dEyGWLAELSseYbVMwRBJkRWsSn
sN3jSgPKp4LT10HbaXH/MTurq1VF2uRJdwkc7ho5IEc0oGx/A3KxNWQ7m2VYZyZh
MQEyWxuVsWUPevMzQZ77wV8I1a8neaOyCkguL5A6pLORPxzuimy8plVKyW1YJAGf
DEsSELI/sdliuksZgrzm0qwK5v4gNsm1PbUrKZeYQ+rVZOmUVoFMIBz4WcY2iBHC
siJ8ZE32KcjjJ2PjvRur9YjhDvGCfgVN/5FXVt3j1kgiEme6JIadUkAvhHEVbEUN
ZCRYVmRr78j9bzhEQFxrRG0jxhJXH5cOc6+wF4l/M7gnOujGsUvvwI26MGwoCqbx
oLn7gW7gv6TrAI1ZERRjCAoq7IEXIfwr/KZVVs3np2qVKRGmtPvSCQQndMQOHV7O
YJ+7EZ+7TIF/GLhgIRMfLFTvgZ6ILYf/LeKxq0XN9Uc/cWOdqW0T+TjnD5DVrIzT
fhMuYDbJMD8SHZuc3zPaGqt8Ly9P4rYDGj17C6Jvfy8RLhsfXXU68VkkikJCL9DX
mEqiJgf8TfUTInsMxqCtIZgotP0Ho/tZpNTF2azAXbjnw/6/pggbbJQASolRAuwQ
OfKwMBZcbkQ2wpymuLM54+eNKr7qjay+LKAClev7J/YuinP40Ditnlc7CU38fJwE
TqZfXjWucn/v0IBphWhzO00u0HPOcwZKGHzSiTzqOk7bQ4BVATeBsqUyX/53ECXy
dYhwF/+6SFnz4flZj3HVU4F58r3PK/xlrKGw56TDkibGapq40uSLQ54aKc+0FAsn
jAvpbHrVrA7MHuiZ7P0SyXaIfzsJQi0J7vQdzzQphTBvejmrTXlysTXMhsex3++x
CUTBhBs+lbDcDDR5wHTSA+AG5WYwoAHLO6sF4hHgGGUaDmHNq/QEqg960bo9zQqz
I2+zuqcvNDFjrYycnWF1Rg1pSQoE1OZxAkK9HKzJiRzVBuQs7Xq8wO7ZZ7iRQrlo
qHcdmzb+W/JzxW99mGdleH/fR8WJD6HM1lWnX1PhRYm5ecem+a7uHO4DPvnqc5q0
4rlNIpb2v0Q0DdkY9Z6+wb4uJY9j6CEGx/GMAphzEpuZHR9QMzFg4715qcArTHzj
U15ZiK6S1P92t6Zch/Wg/XjzE+8MoIwrgPN4FCpg/ps0Kn1jSRxzFSo8rNzauyRu
33xiJlOCTW8L5w41QNNidTM8oGSS9rewtYdC0T2+ENvOxVYaJ+cALug/QRTTxn/0
KUbQ9IzNdwabaWZhkW3t5vtbkXT1GZnKwP9fBcTKG3RcM0T2efBb8YAetdExDmaX
y6ogD8BNz2k7P+cbP/QaIaMgBhTMSxS9x3bH+CJwqn30KWKbY2C3f1MLkgQPJbFo
naoQ68lw2WOnIqyko7d6N9nX51cKFZW21Da2Sm87RvHsUCgnOQ5Eb2Q5jbf/nz+5
Ooj434YD4+0r9/o4rqrxySi3yphsrdrAexUoNuvCRpTYHuRnjcLLHYUmej/t4Ig0
hruVxUFy/CufG1JAM6TKugah/5APPa8W6Zx7aaht9/R6ylI2Lex5OlRD+z1v692f
OiN0VHBugRPYciZeeN+BQjrar5C4m5QAoYAWp4fJ4rntMjuwKz7nysO4VTOJIafA
ObIls8LCDhc3IcjdTXAhXJsp7rybJd/mvUHL+POlx3UiUHZRvdMj7mDdNLzEwNEe
GHu8TqWq30b0pGSRJwj/OGj1Iw4cN3Es2H4R1gScoRiLQK1cWnDbIDe+lq2aDzG+
2j2P/40P+9xM9loJPFQdqMZR9dzSudjmiZlSpVVJ1hjwj0GD2a+CMKSL9xih9v8n
N5CItZPEPbrha/hgiTSDIUw5Gycg7ATCYiwfqYI2F11fKHh4iIzu8c/NpZiRj+mk
YVaD+npDyVZ2YbYXSppb/KpoMCL+LfhuToPoRiiffZJ7psjVeQrMkC73SIVvhIYv
BXdFl0x5s7wvWHUWGkRW20hL1ws9FCl5G+fUOrhcWNDOQY3js8/Re2UOf7IPiqRm
aI2184NCjsu8kbT/TsPR55D7wU6d4KraPt7dBPilVQY9QZcjaP8cjokqB34s4pj0
`protect END_PROTECTED
