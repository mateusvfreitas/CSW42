`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+MStL0algbqhaX5o70HUYRf7WlNC5BQByrHJi3utjzpWV52WGwvVrGr+73pt5aoG
ORHyn3ayvMcZza03qaX2ep+zuRQx0rJvwuYWQzg2d9Z3/kJOO2Lupab2gGC7Ba8Y
S/DXsfcW0m7on50VJpDqu6t5s8dp1lQtiuDwmN6jYOhcD5n4603nHtVt7lTrfvzL
+NF/MFKtnxRItZeuT5S3H9YMYCpo+shvuvNq0u0x237dsT5Mz1siO2cEmqV2nFHo
b7OIUNzuYrpQXw3YKVF0BuheIRU6hzhNb7EqNoh3887XKg2O+SK0T+fy4arHBpvE
mEKCQghTae5JdkLr1/Tw3gfZRBuOn1caOCHEFjjdWe2iGkYbXkxofpqMKM9Qj2Lp
Jjx76ur6zZgxzrg5sylL1Z4b05Xlv4q5qLRkc1sNTsU4TC9o3IOLYqi4mFZxgxyG
hef4xdJXsB7vMVozmBDbsxGCsRu44F0lYNgKvUVaHN5315t1KNGgPIcZfrknDdVg
hN7t1ctH+Nm3ZB2b9fou/y31xoD1ZhhsVp0fF2BWtpA16XAdPVUl17Qy/UWtDe3o
wEaI40MZFNBUsIOUzpRd5tQBJXo+iWz/P7jWesV7gTBR6/lwQT+BXyzPwgOuoVSk
jpIOS7he3AfxrRw+5yBSjDhEAk7irRL+puBxU/93GpGx1PV5XdDl30wRtbwTUcmv
qHUzNf0Y4Nf+ieA2NN6957v+bObs6Ev8FahP0xkdWAW0f9yy65WVgVbjET7HY1nI
sThb3tJAo3Sw87vOYmZfL0CUSPdJGI6gaIEDlsR0Y6iuQC41dy7kR8rAS7dDvw7M
+mEmItWZ9AB657a6fViBpp3Swxh1zz2uwpRcXN5Iw/MiIXd3ddk5EszGSqZXxQLh
87Se9OeihD5F/8sTOOY4rpAiA4I1w9hvUJCEEovAHXpXUTDIt7RCNLud0XzhxN8U
qMs7yAA2ES6A43DG3zPceKr/2tSvKofuX7i6JXyR2GGT5+62QE2VqNy5v5MUrITL
ujrhRay2ST5yy0Nyx98KbaH1ZHxX+JVF6ZaHk4pbKpp1uztsv1JgCpjcAq4YOfLw
APdHRQrnVhExoEZekwph5TlBI1uGPKFWKaQ9FKCec8ZLPFnBQevtCFX7VEvszru5
3FqT6F4GP1DJ6KSTNaUnP4MunFV9mx/P6whNuopRPjjQwiZrUQULBXlYvSQbx/2U
GH+GAqHFf43s8L5Qn/3j6XA7XsUTAZNmVITqtv77trbjGebijzy8UP7DMnG6BqZL
H4JHD3NdcQ3nR0dW/1fJM7l0By5+vR6N+9szBEFCbufoK3djWBfUoCjH/yj57dj8
rGcuqC5TQIlJmrJ24U0MFuaIvKd5N8TOfHBDfOGsolkFpmnw30vw6lNxh2DP03HB
ybzdBOO9GQ576O2YasS++kEqYcBJQSEbhshZsqlKkRVB15sPvIbFN94HA9APhYBC
jJDXTVJ0Yxh8UqM/cYEaq+Pzw3m55oZsG2hPf5/p5Ur7d4zeOR4sYCIkqlARB/nV
w+jtvI85lEtSE8zCpKlOlFK1iqKVMo1Z0U+hKDY+zWWaEWw8P6JhghLDG08oq4MV
HBhRf3c6ftxmaEbGlhKMGGhaw4i2siyH6Az+xst3qMsnZ21fSaa0Z4H6VHUNUe1+
C/BSDwlx6rJfuALKt3z3oqgGhDhPlc9iYUs2rhSJHRfBB6zqlLgG38LxWRIhE4GQ
pdeAr2XzfO68f9BRWAmllnv5AYn9aXorh45D26ZGNuebdJqRpj1qcId5Hukg8syL
Fgn64wOaQk5CRYWU9y5GLiPQRFGc1YFsjl0qiGT0RA9BI0QtHGkr2dKrR9KFaxY/
0hIjIxWo8v9sWtF2CA5wsDHrfyRC5oPz8Mw2KyzF9rE39jloj+dLyfPiz6UDvM6m
zpIICq6D0oi7FncS7SN9u+VTuGct7pC+pGoJB/U+hobjgPlAS8C+opJcQoa4x8oB
mbTjJxmlLzsrUkEcxCXqVVuNVD3Ji+NWniYnFVwqfcnmwsaWj+1wV5nynjIdR4nD
tvOo4yiKNwcdc6d43+GM0mF7K/1rJ5JbD5LkLCJnb2hgbb5rEbLOHIxxJnBSF8q5
deO5xbShh1YdfbbHPI4qYDrUx/z0MHGV/UO3zhvrsqEVZ50KYp1he8qupzzL1y3c
TrPY8h1RJHS9s7KCZMEfKPtYWHpjCSkOQ5wEGRrIy7kBiByzZt7e8G/Du+VEqf+u
ugzP3GEUeYte77lpfyoNitFMPdUGtibSAEf/5+0x/TGwFlmsNsBXBouVe7QQQ28W
8cn0dE6cA7f3PlM0mjDMzbixg8dhp6UHknxj48EqmyAgX1SaJQQ6++P0O7YXWzZM
A0K7v86950gR8S+++pF5eFz4wGjue40Cn02YxjDEKrMywNv77XG90pyNdJWDW4dR
UA1OPQxe0rZm8yFaIoPIYEO6PHFRKLPVBFAneuKp0PcIQklYdH9Y5DbwcTVcM/cA
IgNPHDvqugRnQrRUmc4iEG9i8bldFtGv1ze2MaLTvO6ikVyNYxotkUWX/LiRX0qS
fdGJ8EbIe3xwFd5qz4BCRh9dijEo4zQBpqtRenfAov/MRFixX/XUZLFt8pSSWciq
RUVBukGxq/KOvOESxF+62ltbd7WeAtTmXqXLAZXj2yB5LoqMcnraoAnx3/sv6Zse
WjniCmdan+mtQ3Tpahe3mCcF9Ip1DogUTcrM0AmUDDNMU0wYCN1kAB6/3Taw7E7B
/KEpJPf4y26GlGojLwcGESDW35u2UL368OJ8tLnbNq8q8bIMmtziLhr5Tif/2hoE
sPK5nubqB2WVDDF9UOV9taqj2ne5x+Uh2k7c/8WzX80JzxSlanPC/0uHipVAz9rZ
Nf8H9U3ZduMV7azryIP9bYcK9SU9dPmq9PM1BACvb9DsD1pKU1TnWfsUt0wBvjVr
3khhS7yAunJScpCGuejDpv66NjqWz7/XV8JQJN67KWRLR+VklqGT7oYDp4LliA69
EVJU2Coj58ugheS+FM9NaBeYOeHni4oEX5uJ/B0UDQfBT2qPcNKdGn7veWo1QLYz
QkWJ1vouTzFQ8bXI3jHr4cZ3OYoBpTMXBaOMBBcqcRKsoJ4KiDxTqMDRzJ9cpKia
9J5BKNrt6cWXKSCCMoAUZoPDwa35EkhK7RlYHTb/DY/YVMf6xuIVISh5SIuDxOdO
+yZpMNjSxKn94paDOexfY0Wbf6zm8dAGTe9/K0+DJvbLXW3jZuGE222gsJQsFnkY
+KYRzPBJzyV5CBFYCRhYYndxzKCUiy+lzMN6hy1l2QFYtYjoLwtZLosfAN73m8Rg
oQf3fZLDEVu+Py0yu2jW1QPsg94LbdJaLPZM2bzt/8pjZvCt0ghHeQSOVfOxyK3s
YWhbCVumOiQmBB5Mb9emtSsIIkzz983ocOTnkj+RDNKEy3WRWKYSHTbsmsrRjYpX
XbhTCTLfZozr1+s/+TOGVnvQ1flAWvneUa58JxHvC7mS/P9eig0PCxK8jnzxfQZQ
qkRkmEdvW1WNUOAO1efxCOtJUeniJoSI6UpVQz366pnSK+CkmR9EhMdfWU9vTzPA
uHdhPzqixPpj17nWbD0vkJ3DnTSTvH9UIQRKqgplQEpufrj5f41zX51QdRzlHwpJ
fXfINJ2xCUEcsIrsqLkfc36X/PCceGgv/Uuwj2STvfQOxPCxXjCh/4CE5OzpfpoB
I0AjrPCm1dPmsXiERdIa0ygexauUd0hklJp83N67yihEwuqRo6/AZl4XzRP2sv+F
LXGvSjTIxQg3UG/fRURU3KngLhiXs4ym7lRofZxLSLPaO6ES9kTkt1J3NR4kwy68
2l1UzWxaJ+nedgnIaEUbYKpAGuFFxQNapf5p8kWlpnVEVnOR635Q/t4MfxHoGkf+
U+SBdeN1rGwYbg4yu0upLHuFQ65iYjDPL6q0hQlhFZVCgPpMauxmEtxu9qz9YVYg
pvHI1lqCaIkpeCAK5bx2YN1ZSI0mRYVZiTXt9Nt1uzTxTM8Q+NIqlhBRmbELGrRw
RdcWhxe5uFpa31Xy24sewKiqnrT0Ui6uo0GJH1qTJ3hTCj3jyj/mmpPEhQZbxegb
axtl9H/p+z9sCypzdaRpPN2aGSI7VgrZc2qvdU4gIRFUcS/eMEHvZRjl195GF6pn
PlEzaYHCANEm2B79SxsT4Fejpb+TMvUP5iuzcNvdrsAU1PFVP/cE2PjWlf4xb+YZ
rv6AFzTbqFwMsAm7BghxPyaH40ZnoIz4YObPve9j4MNE+n0s9Sc1CPu3N5PtUGQS
O/niHQPN3K5YpcGPtfOGk2WARuAne9ZJnP9J+LzkkxwBWecroILY1MdprjITu0Vv
FK7gxPw8zKH0FVlazg4o9tOG9Pz7NxPGYISO0Aw2aDD81f3KAx0JO+tGJGSs1ERs
M255ZXziyaHtI/UmdxYuino/vsgRQIziLWT0KWxGjKyww6phbezeQQVFMB5WeF6o
n5JvB5u5MbCHg//dIt1mCmRfO2aXnEteFuEgcrVjNiVFcWOP5K96hewp3p393ODD
BLehgwylgPsUdv1KrKTzfke5eWawA4Z1VvB98aVwRbs12bpZR1a5Ugk4YAs/yXL2
G+Nj5fByCq1XyZQD9fUUVdb3IBpXfmpiYq095IqWGwXcL9ZcIKra1anjSPZK+Ko+
U5Ml2tYXZPGRazjKh6P1BYN0r7XTeUquVWlRhrwwdGXh1D7N69F5VJXN7WWLa/QJ
g7R1MHEG4rkw4BYpY/FHnu08qlpxKmFAmlELPbmZ8AIceido6djoKUjJK1JpVdq2
H4rmsvkCmwXw2pBR5h83iVHaYbllbVs6wHmHaRQxx8e8fhcxsGxeest625rENCFc
fx44XclF7aWw+8e8d9YT0+3/2Xq4wYBQnI7hBNtZmQ9tlxW2Q0Dh5u4lkvpGEbpe
uiM6zNEkQwipzKSv5tTmPfgaS/87Q5z1gUApbiGjjgmD4/1CJzPcACCBth4ntOAk
tMN13OfpJD0UQD/9XlHjBXcCAg+SJXSmYF0Aih70CSB7k0tyIQRPSudzmNbdM6Xh
P0nOs3su0kmLXzkpfcqs3HZeJ4LLQ5oUcLiLMyMpxp8kmXPdpCqTnv6btDIo0Sq+
m2JodxHlnDfCZMxUySTh3k8S71VJtbmfUE7/anrdMkhmNlPtHxjaBklZsktc8cug
NwB281kHlFolyWAYb5+9K8Tfx0xbgbqbf8zw0fW1IeImyfeiYHos1B/IM3LOjwHS
y4rS3zHozhdcLOiAjuW4rY3UIXW9CGyRTmWu6MG60yHfBbcS5fuCjmvadfdVHj0w
LBEMjqPLqnVcuZzSNGKd9epN4tUrcxbCe75BJZPHqOD7DmmhDL8UaNAxUEHINU//
/49BXeqE3I8aHU7U+BI9peADYjvV6afymwZ4xxYsdbaQsS8apUb63MYJbqZSCHuA
m94LvwjOKU8aVpOdWuq4qbkHI6u3dE8BAR9CMHKBYqW02VhIYE1KqE0vpjecmnX9
uzrzaG2liKXmvoOmDu6Z0Pt2inbGLY72mIE0pfLxxSmcrU2TAcmXzeYh79u8SC/b
0nYVCZmAHpZOqPciXEJs47huRhYJow3Cq2LSTbKIE0zz40L+/cb7B2i41k2/qvNd
pGAThDacO0eZMqoQb3mWn/Rfod4JhAv8ighETg7RcIp4YB3tlpIl/Lro8eVloV4j
PBGIRBu1n2/uuKWvYerlo5pFXZdzfJEPyA933y7EmImlse2hpMVae3lvg36hj+VO
B6gHnVKAakCKfM7+3YkXU59RuptynOVZU+CMByTPsnsBV9b8imt5arJ8vJj2rd0x
mifbM8ExFCFHWpal/rvtOhd6Xv4WVMnlPobMxGj03rZxprCvSIbEroacHJd8LhQO
O4uWB+/O0pWoan3iGbZRdQNMhy9R9iwhm+3FtRK96940SJu/aJodEZ8X51+KrkWD
1lM9LRvSj20KwVJ7BJy1HanXm6JmiDJS0OGEX3OFA723EnfWHTEach8zaDQhnRRX
lNq4PSQK1HIr3c0graK3K4KWSl2scaAgRmgc+F6rENM=
`protect END_PROTECTED
