`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2Xl1vz9he9K1tQJEwWOy4YVS60wjSXyi929N/rRU7kDIF6CBajR6omJvyz7guTQl
FpM6SfTr3+kiC9p0XOzV8IwoOQgypTYmt4oELFMGKuvoiAsgVcWo9pdDV3aWvvcf
cYjcrMXH1CL/VFYnviNr2Om7hGfeJfaxAa9JvqyzDl7O+vxpWNdHQ6hd5EopnzZv
S+1B8r5ZA5fOwPgTTuFPq/IymUXZidokwd9VTw5+fd3mclSkKbbqHhpry8Tm/vTu
Exw6HgrrCgwqmGnxbq6TRHSAnIbgKPrJRQ06+bXgsYG5mqYVdJ1bV+MU09P37oom
LMZkkoUz+o+4EXK220Nm/RT46R00eck6WFNhiXNfVQwYBkS9WQF5odB0qWimh82P
rbZOD85nDbDeRn7ZYmqaJ6bsSooGiwTX2rV9Rm7vyim+7heyWbGkakN3Dcn7Zbxs
oPwp2AmKLR20OPY1r2H785suS0XrQBYaeIIfq2495hr0iJjTNvlClgmlZzTwK6mS
sAyhbxtz+q0PjUwpJ5JOtrMw5tP3hAWC2sQmiS5bFFYqbIq9JaGLBNTNJNM7LRej
mEq2SnY3roSyHeia6Y8EIqdlqiuo1BnZq450ALsrsNfjDH8asbM/mNWDDTMC9/ic
YivQI6qkt9BqGuOBo2DhvLZi/sDObezR72tJ4nhBnA25luQldj4VYvliUv0vKBYi
lfwRCtXqIDZ5sOSOrah5asvJTIavoMxkWD0ECqSwqD57fEeH4qzJARddOgwWutLa
nInxspDcxAkvrjuv4zPMFmDYg/rgMJ3zrB3P28+T5mO9l4R+1vKUN+w4MQkB4zxT
T6njJo/1j+r/uJk5zdZ6HOecciBrhRB+IQLkt5i49P6Vh0eR7g36QTWRUxjzLwmQ
Lb6pgYe3xURq0nYbfl/E4yVJJOyIdxAhaeYijU+AMZbqVBAtLizM5KopXkfS0v4o
vYPmKaSIWPfaSJXcoWed4jBQAydNxB1R/UTf1B+pTG0a4tzTsm1eJcc7co9rrKub
39XADFQDhd3oSBmoT6mSHgROfjl5hEvvsn/7wk4Ddua1c8NMMO/rzLGipqTVXCMN
2/k3b+frtLD6FQyQAg1BiZzf2S1Yl4yhKKPp9suq83r9DWU8iT/P8wHMfqDXJHo0
UbGbLvRE5b7vH42Ss34O4xRpQ6EYLHWeZmyvxm/fdCz3IEJwpgQmSv7JCjCz8Ece
PkmKN3+oG5h77bau/DCj+EbdyuD4r23LwBzbHt1FrVZTgP4chDnenIm4nIKiu86c
6358MxiPjF/uNZ3xhR+NF8264XeiyOKj7IhJhTAZ30u68D34FVSJYmpdSviANK9f
15ZPKTY6lMXQ2E8vKBb60GgmeE9LE7d49WCcPxgQqnu7R2jhdN1CmfO+V0f2XLaQ
Db47s6QaHCk4erUTo3/NMc/Ka17FnjPlLTBMhE7mvaLDz3deODsTQQr9td9kW3Vz
Ws3nOgCXMrHqGbGJfLrwJ8eVCpB7gFCDkg1b4rLhxT/ItmA8tY6PsVVu0idJkohU
e4dOmQeatO4bEJ6jjfR9wHzlaJXU1eb38dIcrgY8NobB7zjh5oQCT8gL6kGWoTX4
5Z7od5pXcQxVcrLNqc15Xw2ThfDtJ7aJTp3tarz1+Pmq29O0ElCeeR6rCQYYLABJ
mIUAknQsomZ35/hU14BNtwS6BS92p7HXcaPmYBpNifjs3EwCt5Xe2Y2wjAHM4wgG
mumB04wrroVkbiQ8l2lTpFDXC4docVa27RvG25f58WNG9mFcVohx/PFTO772JjP+
1qWQYSoWM/8cAHxv+6SdE4fGCJKleid4no/+NZcpNGR09eGfGcXqM61c7Zc+1jFh
TbTF9aOXCJIKRHQZeYxEZiCzhTuNua5ugdj9A8VUpL1OUPG4NpjutMNl8rWIkwJr
pCb90gNNO6CyugTvOZhMC3ZcILoh395r5IVZACwsMOl5ehbCb/Ybjd60/g8PX0N7
9fDYvAkJP8CofjS8RAQFPw6lHYCvbQpcNU8tHuEvKsJ3yY7SdzzGmHpIjd9Hq3nn
OQabht5s6keUNWSTjNjeC4jm/YT9+DBlmK8mrAvbAcO+gkWl1PCeIobD5E1Koe14
eIQv9fH1++9LmhTjl/i868YcKLUDXZvMxOOiDr7iNs3blgB8d/7tx5Qn3IlnuSPv
DNwwu4EDLSdwHIzbPzuZQ0XCer1bhLp2k1gF2kT7tefsluK5WSgHTsraPW3yYFzG
qg7/TVoqyFmheaWEhqgWMUHgW7C1Y417ZGnq1SHHoQlQVZ9YUN7Ppl1gCNFf4rE8
ebJgRW/9Vrj394j/ayd4frhS1u+cF0by1qPR3aYpQKvbzK5jsWu5MGn8Cv+tWwQo
X25q0fyq45E3WBSmVx+RwOtcbvgB7f5mr92vG1g10YgubtDbhr23bOnXH3wKNqRW
sLKtKXCyadbKjHLJw+fyLZqOvoFaRk5tUVTt8jYqiGXBD7wf+jCzsAbaPj+fAT2S
p7Q0EPy/3Gx80/Bb1ACn4H60mI2uX4qELVcyPB5ZEdTi8XI5Rfqn1B0o3g62IVA1
tTfPVO/l7fi1kxM344qVMRBYlvpWV4KnJH5cafOc3Xk49MEmG34RvOiE0EEr8IkL
xJchb5KSJFAzG2n/dyFXBOaCagsEAl678lFWZDIFHWPxW4oct4c1vNCqlCxDPTUC
hhkM9likldSlNYj2g5OB45QPU0puYSgVbEvgkC/tjN3lUEArSLN786sbd+3Nqcun
tnyTA3H9cH2Fsj1Yf99j9KZQDOD04iS3zUAlSkQzVMxVgmctTb07eHJ0LPAN4FvW
T/Jq9jUK4zWMGVOw70KrcmXf1S+v/r9xx0RXjeNx3n6IfEh8UVcsYdLDym9zWsbx
dk92g5CFnd3IjXniF7VQ3J5Tw2acsMX0J8AgGvmXDS+VkqWzIoNFPff3fI7kaUgr
3gWdJt/T5Fd0Qw7s+3eBnqiCKpy3ADVRJWN2ZzJViAfEcgCmtini2f8d3+NmYxIz
Lorl3LdSynNjyo17rPjtGMt41Tcc+7JCUafCPRNAkQXiw61CinoddIFjLOBAW1x0
yLOrzWO+Z9dRn17R0bfjnKvT/r+bNgqF6ZunmpD4O4w3XZYNS0OrixKcnV1N4KTr
w3sYA1RPvpMLo9uiPTjSYv6yACyJbCIFp3NRuSk1smz2Yx6EcNdEjJtR06bASNnK
sHPGddbwbngU08PD5kSEKzFFTBsPt17CIiLrJLL5n6ciOwhK37NpMV8lai6+tTOB
bpw6MuAhJW13u82YbjG165badILfh417bHsdYB5L0GL2TE2OkMFUz0vIpB+o9jxT
7hF6tC59fCyjCKwIclWD0qf/Nr8N/ZL4lK2OS+gsCZSqbp6rGtebATv4XCckVZZr
MwpY2LoSINEjmc+pj7vTmK6Hp3Jhhjj76qHFar5QLWlvDVkbhiaMdkuaC0zWX2eW
O5RX7GTiEEEA0njcu0EY/UHMbBqI6r9bUeWhGhKOmjVEXStEFz9cFmimgL4Th+14
pv7eHo2Y9vIwbxBGi8U4JMABTQ0+Nki5Upgi3A4Sk51gV7KsKj+sYOxHby/aHTDJ
SRdrRjnGUVvNarLYKgouVjp0ST1ScfhyeaOcI2IU1flh4QyeH9PCurl4eaqUxFSY
P+q1FJoiJnACK105N137MK6O8x5Cip4ZMDqjJoxCe/QiUGCWOuzIqRWOMDwiBpnw
/rqKrHYVwfH1PXH7BExzEZGS2ZjEpYth7NFKBSUzXLkcqsWZ3F24gAaHRw7OUpOY
0qQAn/Y0tRmn7w0biRJQISS8Ifn9tEOpE0ftnnCUzfTwnWxEyY1GNIrhkpLavjVg
3ACEmANkQ5VEUhg2a6abNDcx1kk378/pCvkeo+ICThK3zKXIPLcl8Le8/1xN63sX
TidF/ps4GH5ZhYXuWiUvO2azuUU2MOt+9+kTmmcCoZa9EVBwjBS/4UCMUeZk1ysN
jxSqe4utV8jekfrZ9/FShuJkFCaIkh8xBQ44csQqfcnyqZ7i1bb8qRnrenZNv8+L
HCPKHnN5sNXjLH/CG69Xo1/9ohlMHyf5vWMmY0JDOyVH33xjs044ZsmQXlwYOhE4
FQb+4stbay6nrzk+jthpmeh/ECrN2RvUVo3dqp11Gzaq/kB8BPqXXQJnzxuPTvLu
Z8ndbwPR9vw16VLPGoFwOVVcqNzyZr9dNNgg0xl2EiaOonRl4jocuwiTZoEGOf6o
Wcv2OXbmHXo4N8xvvrKqn7Om9XKLzFdsdJzaZ/NSWwHPAs/TpSXVcFWlSZPGmuHM
+57MzFZKHPe4X68FteSPHu/jCfaMWRlbSIVjfQC1RH5e6pH96GWa4F83yeae8aWc
qn+PCtJqPFJGRvcFfjZoq9pFvlidFqwYbEQAHB6lK9WVdrAhyMDnxbmjm6pwdglz
rW/cLCoW85u2/0Zl7mw73Ey2MhW8DCWqnY1kdjcfnMQVx9AIrGIBnGPk6YNUSonl
HxXAf2ddOSnUjijI4WEGmwqhfFmANQAtaVqbHW4hpnQ/DGYrd6VtgqHCFzJ3Kcfu
rbVbEywJM2MVh1ir//eI6+Cvb0qlBn1XWciYiy8dj0Z+R5d8SzDs16a0ZJHJqack
Ka9j7hg/X9VXZDclV7daQCWwpcA+sP7WXsSrbKPhh+rJrgmp/cQUwOsPXf7S7DMi
guGPUKWnUCvta0XxOfKVf6Jksc+ATdFAC6bbROc8pcKBGgkn1UnzibQUKR6MC+yi
Hot+O25giY56CRLBYv4LbEBpzaBtEVnSw+AeqnUNLJYA4iZd7WfjowHbtbqCh5Qh
OmWC+8Y5lD7l7C2rZSM8eL4PsPQmI7XJft079qhxEKe9sPrkY5WVxfcJygzpGxXC
bafMSA2grDlCPwigJgoUqNp5KA+Ybo9fmeuPPeaOQyJasJ+clVo1Cb4inSTlAI8B
2B1jCbqsMYU23ePuBJGxluCF02yC5JAs1GBRAFBSDzJx5s8ttf7Py3TzZ25ItTaa
ksTdVJ3MEHI4OX8dnitE82X7yHWc/o1oxZqNnoJxWGXlhq8o4NezOUNvRcdWa1DS
QexYawFYDWd4zB7FUkl+CZcJGGhMKb22Ezgnq/B2cZTnjeClgDRsxi9cGQcniGuB
gNq6CfKhF4CLZ9y/KaygO6eOCxUj5liFT0kZuUE3NrgDfCyeisPWqzYbdLgq6a2H
h2klfN3eTQF+zLxh9hcFMyruzphmod+ZvtOjIYHVK1y4mUvCB4HlMwnImw9+T9qd
7izMoCxYOzgHvB/il8JDy2X3jdvZD/ltoFEBvZonIvtMzHgMZExvlTNFgaC3oxZR
0mVvH9RedPKoLbApEtgk32G4BG3KxugJ843UMopmqgj8iH30mNs5QqBUKX169lZ5
XqX7e7frqCn6glpyAmSZII5NStGsVYV6QUYGonKsM/vydhg77rE2TDLqvxeUaXVR
fdYW4Se7Bh+WpHOoZs7aHq+B0A5X2Kl+TUQQcPpoI9aLPIFOpry7NVy8ba1Yp5IF
pRrQHxgnUfauIaJfgXbcJTQ7ZAbJb5/VhrK2vyAu3jS6J4sykE43tiPob1YFa28c
2PvKlwhi2av6yllkD7lj4Lqyj671RtJDAz3BwG0/2QqmliE0inqf/2G8OxW1paFX
pOalJo8hGIQPgieoXJX2IiPgwcPf/o2IVSbOrTM41X33HGq8PgLzpBpmu2K/HG4w
+otN+JIef91/EnJGD66HVDfcYtpvJ2E0/qdhyrpA/umGJ6qwHiIrm6Zb+sDxbXLA
3jj9aQ4Yt4B0vnVw4MD+Wx7enFTht7rRSa+J/iD3DuCDsj0MynlYml31FD4kHIk+
ffo5nbaw6bc4NS7YyIm6B7tqSx6oa4Kvd1mKk4vk68ddJ2o2zRfkBVT7efvrNnXo
VdYr200ZUQuG6OmT6QHxlPM4DEQL2mkx13P9txa9hWXxaNtUAAa0lN7uOLPWa7X1
hc0eB7igUFMdvPUG5RG7bcOn2kY0yAWOynVqee6XxzRyXPxI+fCwwEJmtQ2lsY1w
7TTx5daX2taoVpOIiCFM56UXXkf4ffLRDNiMzBLn/BnNcVX6nkeSWCILPGCtavE/
bQm/BQVeXpHShE2BAWqg0k/bMbx2IYFWQ6EPHQUbB3NSG/hhZytnGAwiWpaX3TKB
ta4669ggfS2WIHDmUvPBviArjNv1cRUnAfP+IYC68N3YW+aRj0EhQVH85m9GmBek
Q37t00uWTBiKh/U413sldf8yLO2GFZhIsr26XOvUAJwBbME5dRuDP52ftGKr74Hh
rRksRSrWNSQ2cVzl3kzRmLELFZn4qfsg9dPi0fB9haRaVZg6b8MUWTGJCN1Xj3fH
isLjvlgbSjWukl92k7yL5ClG7TczUytqHKRCd79w7Km3aROa9uKXTyJ4FyHBq7EK
C/CFG/YHrrREepXjHK7oDJSpmRXdtdpua+NN0FRq/yUNSWhOntjIS8jrzCQMhVWb
KOCXHf7hvRSlc5vXGtaH7gzEjC/WnW1+hCAj9guxzanZWd0sV4LgL2HVbjJ1jzK6
M91g2hPddYHkfNxJE0VWRUCpl+w8lPRRiXnB7dTy31wEV4kFWEO0vL1mCyD3xuOx
w7V0Bwuv9wMWO6xHuQ01KDSamlVeeUYVUJ+mVMfgdmvk+WM+3lZY4wpkBztTQ/q7
1UgQw76vfKD5Oh5Hvp/m0ghN6uGUVy5U/9jsPZza9ro=
`protect END_PROTECTED
