`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
1YF6cLKeRAlL5INhy6DCg+4Z9714SfOnHw4XQOxX6YkStBmVDT9EalEMIGP0XlxL
QZ+KDtoEZ3LV1lEJ7s7J5RojHvoToHrMN8+Ah2iKgLDSJD/z6+R8boFPEmYZ7VuL
boCFBUEDjYcIWkO8x+DPlxwnDko/ayTIxPG38Vsb0O47YdTBsaZXR+N6CTdd5ko8
4dEXxh9s/H3NaGxgqWdFrcO5nfhiuvXhixJtOT0mmY6OT3x96c99EIQIlkMAcf+A
EVGeaDlgPtHDZiR1bgiu7qAblhZwZyDtLuyq2EvAHf8ssLBTSfbQEErw4+N7k3Q9
lRUacTNN6i5hML50/aPIVOsYXrH8Y410PFHMM4YsXOyc6wCIVL+uxnHYbk22IbHO
olXqJH3oXqEEFHJmBTkNfeZ+rUr56fhD86dvcHaQWPZJuUZIDiNRec9NldyN4eo3
RFZHk6J3sVhR2Ya8CrUYxEqiEB0nPOpBq9vILrF6nS5/+TUzZKQX5LhQqT8y5I5K
UVHIA9D0kvPXh1aItrpftQ0wXhoiYXkEiznbfovaBBtGue0acQmCgW6U43WtRDuv
EONSKKQuf/iTpQKHVrLewdp5zIppWB/w6eUIaZkIzGqHohCY/4gcB09RG0tcVNHP
TyBX//NOHcAKx3yr4ovzLszR4LTcRYW76ryFol2upkWYO3jlDzjEUp6tgWZNoMN4
ff6cwqVEzRwVBekI/9QqvzdIGwvz2F/ELH5DPU6OP4IgJJf50yULdju+ASG4TDYR
hMckwvNvIm0d7x+Ur4zX3AywXGxFrX7S/GuOtb5EO8T85ORvLlYP1Piuv/1Q0jdz
Bm6uxPlUC7C92oH1/df528u4cjkWctPUSBta1bd0tL5WKoPinHn6TdjA458u38Uj
yWut+QBE3sBzpznBtWhB1zgwn5ZtVqd7FonN74JGmkfpLiQTpbcZMaiibeXXtmX7
u/YKg4TA0nHCOA2qAtuoRemhTm4bCJKbPN3D9jzfsarGiMjT4EnkjFC5JRoVAEFY
9Spsdn2VjXDM9pE6QFSiVBFjJCF3EttC8XCOcJUJegwXo/F6NpW19iNtDMuu+TLU
CTm55bAgyyH3ghPOfRy1nbNAG0P+Ke6Xg1Au1xiwSXAJbPzl5TmM9OsSsMV28UiT
L4OGZg/k4uRdUbsKbCBxSRoDR8N+0FWZKz4TM5l9cJbpNrawLl30KdBW2/X+zAGK
cwj6qBnqhqmyFJ+dU1lHb5ReedJr8II5wFOPXye/MeTFqVU82qc36JkLH8NuGPP+
sb9Q6Wdl2EFXEB3ifRfVeXc/MNM6pXgypp6biFMo1tjC4lQ/hCGYZwcUwVnVs5cV
ml2Z7g6Lty5T3aFlKs0ZqWu5dOiYlOaeQePUjkVG8g/IbNcKODSJj5LN5WV3E/ft
mWcv+xkqW/s4hdDKQtQn4bDdJb5alKrGeY8fYHQtKqx3mcfthdaUA9QEL9IJXUxt
0OYdi58Zu3xYcYNnMLHpZHrvAoXEsEs30PlQnA1m+D2Gax2ctdOjNNVkRg3S15eq
Id7GK/qRPeeyoEwD+czMnIqils2PdBfyBqCKRIj+aiSiEkQML+z6lIbdTz9EjZ2r
+W7IzWbrh1fc6ZvMtfAJqyHlt9GAPczT0/XBKIJD8UG78loZiw04xrdxg2iJ6cxs
wyp3v6ltzsVVX6OE0e5w6nUDeFTccaGhrrxR/y1nipLTRtv9mKRWhXe0K3U5YSC1
SMuICB28gfOmq4pqyCSYbqwJrMzllDsMiyRI4y5hUWnwv3K7h3BD5mgRsyeyZ79g
dH3vcvglXtQ+cKp60lCVC+AvesWJpR9WBIncGK/jhKku/ZgqXSgHmRnp9Dm6DncP
g+f+Fp2itk+WCbnjkvhe9of5IREZGwaTtUMg/AFmP+3YQMX/KUjsHi2v5aSFzU2M
HkHPc/eo8+fm7sB7tMO4fjUpYpBnCZZwUgzOUVikbebu1hXP1mSceMJH55vfBuaC
PMXwFCOoGz19SQIXVDIrXuMECCnAfkXmNmVTTzTTi+lVMjU/9ywb5yOg1CHfRxfT
8hXKp+/u+9iDe3L8n3nXCaKGipmr5GAuqT6tQ38/H8tk7MBJNQhenhATH9Ul10bK
mdEHdZersqDIhe/aDLVB3kNFywe6S9RP6h+6xg1KRXskuwRmfuj25OMLbXTTEhSW
Ed35wQSeE3WNIHMqoGzxb7Wjz3BVBlu/LUFihpDpq6htHzR8fq0fZ6BdsymQ89fS
NDdnwNMaIupM4d+R6UZc+I8KdODkv/cHa315rWNbqcHnb5IqnRp4cp8iva/qlLaI
kODpPTzDTnEv1f6Szg5l+GQel3lXt98y4CMmU2CIGzGixvmHq/F7wjkouOwYdaBf
UyW5jI2Ao+b4IiE++xYrbNz1CNnxQejVXCXEYaIdLD21qR4uby5cCqXOzM6ZgoGA
5xapSAoSgWU2GbPZMfZnzob1Hkp0+83YdNpwKByOCmfqg3Vc0u7+UGmhgZjLxm2X
ll1Vntm8/8DAPHtxQzJe00VGkJsjgw6KuVv3Q+h8AZGBA0dwNOIgra13BTWo4oH0
lCPqUGH4wB6uPncryza6MixlFTif6VVjq8eAVqclCurtphfHyGJqN5HynxuNjwFo
TEYb/LdIWuMAGqnQYU7rlAk20MPj62JwZSMcLSMztgDmHfS5tfSU2BL3I4xIniUo
QnlTLHhREyGPhmrcidQpvN/afyRfao47jKAnUw2jiVlW/2Cj9Lz4ddRBopImIcFD
BxphjqHT08ZZTX2jEvu7kFQIcK8VIFAW11CPg0hDWi/beqnpaH5cCRzoDw2EgY4T
D1/wcJ6jocygaXdgiwfth1nUf0KS8ywmNZ6yN+0oAJx5phlmoYktp5ajwYvz8W/k
kMXMxXZZAao/LZLS43GeHynnB/7LpcIOMpAvvVn071YrLl8TM3mON8aeO4Atm6b7
pl10I25uhuxdRNMINwW3X1kgzBz5yHuj8vnIcX5fuymeL0J7uRk7DBXbfIpa9jAN
Eo2RS0lsXKyD4OChk1CTny16lBaRU4qj4b1ySmOcCYxdaGU6fLLXgqnVA/jE201B
NDQswohk20AYGxRi1wjYsxteOceikqDBAgswyqBvuGIBtajcaFOiRaFUd1BahvBc
PdRm7lNAmSMDHgNHxINSgYfz0UqL0Z9T+RUsc9pGnJUCO7Ib/ijbi8AUEAVs9gh6
dA71VoZ1i4+5GUvmwna8pMK6xBFvdc2wcDYdDACy9KTzEVZgwfjuP2D2jIQ5nPNv
EWWvmfNxRknUWrDDauGmuSrjEiKctlwDIBWhbXCtrJ1oFVONlMIaOXV4tH2MLKHI
yVQtD/pg4XfE/rwkFGXqWVEAZ6AdDYRF9mg+u/usiw3IqVZax5asN7wspZ8E9Q37
jXka4pb0H61m23olmqcq9dzdJNhsI7ZS7ROcxSUkZOJ15dMil6chG5PaRVpq+hiO
kZSnzAa747s9YhNEQkK4v6kdF03vS47MEWV9mNssXDk5PIuEb80EfY3shfv1BjOL
SIxbOcVa679PIMNlsRHozDJ5eln9oZgs/aeFtwxwiS9w39pAuZXnnBgqZhDmMb9/
/4R7ogvTW2MLJ/e6R5rfOXpDIvxC7XPakQa+WmMyD9yAZ5R8Pan7yrTagbXWneo1
DYq7n4zfNh60GRJuFnE1nCmB2z/GsOiLw3erC64VcM9ha1jfd/Dkqm/346elBGc6
TRlTx9qDy7D9LEk9UpaCBS9iRDByS3BAR/wvSTne/VKxDrKKz/szmiheRzjJ+dDY
70eo2zXPo2TA1exNmyKXYbgsnvDYXarn5TPx/q7kFuOif1pTWZ/xDYkLam3i5GKt
Di65CkABfM/cwr630uDPxqOvoF60QIzz3+ql2S7G3aUPf6/S8vBhLE2txf1iIq21
G5eklfMJtMrFgrBaXdnd9MuKOougGhdHIjg2YZ/lgelezETu6Tc6QqBeyYkZcBy/
c3iAjqUPegXqNdcqYLnzLCcDx4Pn0DFoISxkrk3Zxq/ZIpnWTzz+VD94EK91k16i
l9fNEBIQhlLrcLoEkZ+IV7Y264U1c7i3TLpIMqIZPzGu/Hzexw8TQVko0LXtwuPe
E+dNsKM/sAtEytdCVVHHFYB3WqyXMCMMZzwVDB00FOk4o6nSRtSUAlaB/C+v2K9c
Q3tLfjCKyQOaqH9UZp65Cd8mjc9cbF4Ax6E8q7EXx0A8+uMaXDoeXmgNa5lhJx++
rdj8vlDm5SOXzBhblNmPE+W0mB8opimDehE6V8/d48rg/0As1kZNvRp/4pmsMisZ
cN9zaNxaxQcPMTATzw4TKz+sb/LYMXZBnWZ+6MJE295KKvkWeeGJb+H2dKqK/Gvb
uOj3eUQJqB3wnDfgWQf4HB5o98RtTUAzeyYZQ4QloG58gQnQzeLNxO2Uh5FoOTZ2
A6/G0t5WMz2VmxPMx9gx3RSu26t/0dpS28DAR6blz8Iri8s2wCfQLpbRQJeG8Xcu
112ZxJRA22/Y98/ybGQUb5hHPBpRP4rSuLqLeH8WU6LtZceW2/WlrPhas461/OzW
mpNbuDquM3XpTJMvHAqNAFHdtFIiC9nrWRxgli9yy6Ts8tfb6PCt6GGP92xuSsx5
L40MBP1ckVNzorrsPdJed4oo7rPtkIEFtcT+yoxrw4VgptglMnHkKacNdUm5LMQt
dXShTN2ojeIpNO9DIwno9/Nt4UYcSp7Fo1okrA1JGKzzRW2uQ1xyvFMXcvumZNvn
pvbQyt/mIogDViduv1N1xlxDcuSFdVhTGWokxCFebnSQQaBucAoO+dZ8Y6DeAMVY
9BG5NYlIZvdWoSxtppqZ2678kP4vjo1nfaDwDTeDKrtc45a52DhwFPVkKviEUem9
SURc8GnrTyJwfv4hcHu8diortlN8VcB71c/TqZvejQpr8651CU56RpCqoxihpQz7
o/1Mk3leIZ6eUargPs1Zan482HvuGMPsOk4/GUSrf7SWVQdaSbtihj/gQYRPfg6t
v+oqOvOyGywg/AsV9Cp1BOqYZA6zM+CdWQxc5uJJaeiOLhCSR57wiRNfR+PF6WqV
tm/wXUyplRNst5Cc9HBXFD+EgG9wAh/TqPudyjN6J150isYKZQnBiU7lY/V0G5Pw
z5KzIX05UIQ0fbWatY5C3x9LP9lNTv0VjKSRlZlF6vld9+sj2Kzgzl5vwOahLSxU
qitTWablvggvueaZgghd9of4zDI5PTLDVaG6recJgGAVIqW19wg2KsjuYmOgyRYb
u/FjAu7oyF1XybG/2+hz3do+N0Zr7Y//WVxNXySRrfPhJxxDNqy2FY2uDyyglPay
qveIZKx5K7SHxXwEe4s0vtJKk2ity16XXX4ZwYu/SLPcihoXgUc92GgsGedOTk86
DBK+ELyOuJW85NkaxmtYvIDfxhzg6AcEzks8QprPCV19Gw4m8bYDJjmCKQLa40bX
oLMJ0gNtaEj2FNJGANICmman1c5J4emU6oma9yCXO5UQckaBz3UHgTxGB902/t8P
NQ+EvdkuLHmaUiNy1DWKij5RC9AZaYaeFWVzd4CiMb4mj5/ggiAN2q+DrCTU4tnP
sLhbJX0FZZ54kM8Q/G3NqmTbtMwPG1185vsDNDpXBxVFBpSt5yPwNa97AaFYX06H
XW6/f4SkYPkVMjqj9gYhYu2LQTTYCv/VLOQyeIIo/ps+8Ot9X39sG6GjqLLOQqeN
yHhehqwkasgg7XmTtPYoUp0V2Zyi/d8DdSx4q0/IMWwnz/5qkSZvjAjzaxUx2vjm
YRYZFmkQ8rDotLnUMuRoCc2Z0q5f3M6swRDLlgDLOeIEZSQeVvITDcEuaefphkY6
tzKtlomnP0a6bXi0gQZVTyhHrShh81V5fLzCzIAQ3X6HSozZDwI+JqGDRer5LdPM
HcEUXqo5m/D1ZEmBxXBforBJRuf9+jLHT763njv2aVxsf+YyhaUqMbAojByc6Pi+
bgrhDnyiXl/rFHKZf/1g54y4qv8vuo6HhBOTKxoZjA2ANeq9uMDcbkCdjwSrRNXo
+HbCHlWiJDP/Zjc7TaPpVUQnQRqdXdZNkWHf2RVrgK4=
`protect END_PROTECTED
