`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
LjhM2ZY6fA2a0rHTeQ12Ipu1Vva/OYoYyIXFkPNodnSBHFDL9LWwKECMFEuVsVnp
lGuSP4OCPvJQoEzdkblSvzLc/2JX6kyNhCSl13hRKw04XC7jSRpdgzZcK/wg15Nk
2wSPfqK00Cqrf6ScEAGC2zALQ01rwlgenY+i8C5rI/8INW5uTDakoDcoyErBCj7G
+TCDbC2pUI0QGHaSqSRBBcxuMNcDxJia2JNPuiQKdQT/1Bt8iV325eypS6K8UfKY
4Twf3u4eEYt0BWtaJb7wP5rEvu0kmMXcAkQ0T5i8kFCu3KokiWPJZeymJNYLcdK2
8S40p1kvuYadSlOeFht8LXCeZes7iPRKWpENm8xlY/kD/huOyQUhAXh4MrTrrLfM
p9SZR/ZuVsW2Wruxmw6Dn+IjefVRcqf25RP0I+SfQBq/NlmnbW/veRx/ZLRkIMsz
3spHm7HXQvkVVxgWWfIpqUpWtVQ+TtjohYoaPlVm6IHwOv9j+OgHaRjtAbGNx3Jf
v1hKc2j1jb0vL2wcyx8o+ESFIoVG95dm8AIWwgxX/wI70QBnhycevngHa0BWw391
rlspZS6MZ6GdQh0k++HluDXRAYA3aKv7rEmrkTCX6CGKt2DLw3UloF9dCQpKshLU
S5G//TBMQdmqSmh2R+dhsEjFuiqMfnh5KLfORtaszcf/QL04JTH89cmSHfivqFE8
u6aIahodeJWh/dniHaUal9rw+twM1gUSwb67rwjkxDjAmPTfvif3QuzeUgONRQZ0
hwQPWzbXudSVxeipDEAl241nyyf3XJ/3r85mHcG+IVXqlSQwWznWT82koIW8kyaz
mNG0xHLqS+chH/U5fHUWL0/j3W9LI0Hct7+rd4PV4kGdnQpCngC/5XAT73S5kf14
hUyFxGMsYER3xA4qF9nILeJ0RWtx4j2hNlzHKn+RZ9iEul9jSpEnNo6arb6CB0zi
w/fsxWvdcHINuSP2ed/FQyyWb98o86jxQNw0J/dxB5Fi21XPyGAJcswgH/bR8tqd
oXXYT5HDP9ru0HS0IA061OonXJN7OQ3HBaE+HoJA6iwIh2GDU6v7pfsJ2IVU4Qse
iBoAEdWpc7k5dDccHGt5uatvFKKPOn796WKeHPlnvTP1YsYlDidt1HJV+J5/bL+V
ti6RXsra7OLkDFXC5G62rNFlKPIncoKq3NxiO6jcegvI2zt2bOrMVL7iXGsqrsrh
SYGVBrpt+h8Y9eKIepYMaQQk7samOvImpHh7QUGTYQWLM8Nz1LkRK7dABLiT1Hep
L+X3W+0WmFGGizaFzxIQ7nkGwp31jFFBKlThgVsMLAvFtaVw6N9VKNldO/8Q+vQG
Ilp9GkxNONye5+xkkgRDZt7X4hyq2jzzu2PmXhjOFb3uSjNEgXKqEIen9KJtxuJE
ab1Rwo8N9eybpxSrRKDjNTJu+UKNvwnbHI1+AeBmy5GDnPBMtgBZYLiskA7QJ5hi
+zhHpTEPjcA+Y8hIrV2gkkceN3tyBxnmcoocPKfX9XkF9ubXHQjqhMwTLojeFgdy
EbqO/0IkWJzOcv9xG3KV9eg9//dKfI1sHL5+F2roLMLAJnm8P0fCLUo88wpVi+N8
7msfYfEzdP19z0yam0jmArPVVw8AdYajj07HMDl3snbyyYZCnIqtadWRk0kqdunK
kA102qSNXTWGnw2MaRD0LDRdu3vqn/Z9jYzk53c851nvpkYcYNbrEgDccdcsFDv9
gWyPcnG/syZEkEtYqW0dLFqNoyMO1hOAY2VXlAB2boY1xpBxdnjf1MflFBaknGPX
SOBhtzl3/XLxtBGRRoQ6ehUIIBLx2mTOKtrGP/F5za9osQub4TghYbk+1g8/GN3d
jKWsbdV0LZLfs3kHGPIiOiq2yj06mR5thdlH6Dh8VQM58jcJkA/2YNd/Ze/yUATv
GkBqB14gdKvRs+XODrqLnW3RvokMIyuKe2DXV08Jt3yWedqxEWTupZhHKcfkuHKs
hvrhWe3vYW1QBCm3LRVSoEooNxVg4JNse2Di7E3no5eScJe+jqS9n4Zv78T9Xsnr
`protect END_PROTECTED
