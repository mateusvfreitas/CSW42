`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
oZa1ox+pipxAzTenlloOaiGm86c5sVHtlmxv5dvFE5ulUGiECe+as+jJ7V7coUpH
FvrC+x55CeK8TkrvOa88/iDYXAUJYezjjpQlmWckBoV4PyTN7ClYGGjfKg8GEYSM
HLLXsTcHQpbSmMoro3KiWAsHTqIyxhKk6hcNV0fnFuAjLv3BFW8Z54tqobBB3sJ+
p2JCLQ5siFFc0QsoD01qCDBSpq3A6LUEwVafQuCtVfb60xFmYzs1WhiStiykzrQA
kUyA1I9p+sWX17zXO5FY7o6l4IFw2sTDoDPYCf/sJmaZHND8kWV2p9k+O7yvRzdh
d40KAog3XBDzamla4DVAkmQBvZedHnexl5fBjibZT4gMuehQnjyi4DcXTbqyKl3+
q+CfQdtJS1PBWuaDW993EbrjkenXg6RyxnnGmb9D+2At8cGrIewzu2TCwgHlXT2O
rQ3eJu9FcHMrHjK4FUewilEOarZhxF1mMrVSQDmdJFmBFkbycsepXHYbMjvCYYMU
S2/RSW9ju1ygKZoZhbtVuxEpOV735Ifs6SkAFc3wiF5xqD8l4ZvrtAQWclmFFrTZ
nreZubvu5OzqH/uaqf3buPR6HesCvVUE/lo8TayEhGcjl1TNwQ89Cjiq9ol2iYAt
atTsVM6OXq/OnT3DlU9+n0ovs5eZ3N0UHFHKNOfa6mZ7wDHQuVEltGNq0mClZj4J
xeQ1ea6CAyhxsxEnqIfSunk6p08PE+l+ntRwkNTzEscFCpQw8300O+95xqbzCfY+
d3G8K74XkVV5estTQtkQJ1SlmGmUYJ5ejXuY0RLRDXC3C9PfLPkfxXc+iaa8VO2/
FozPq0TBI5IQfjcKJPaxkVPfFqq+vok670j/ePWJIM4o/+DwIDGab6pvoU/mYY7y
FYbLhrATXgvfmcIarrSLezh9OGVdedlZ3K+fMK3AYDhXAVmRB50+ELdlYctO0wqf
XNHkE1+C3km0lcbLsak2DZpWbz//JoCnpTUjpdgtGNcK015tTVqxP7R0Wfb8iUY6
hHpo6bKh3x+y0HRovFwKwGCMNoN4pX+VavlZxmL2o/h1DOUDo06JcwpRm7/xukLt
Ts2g0S75aftLI6ZcOgZ/xS6qIF+ywZTm/FImOkK9VLqmO+sbbI58gY3Ybv9nAW3H
PamJAdI9kD1FJaX6jGI8PjI1NntzpyUxx2Se7/bg9uyC7grxiQL5E/dD/Jgi6Hzp
0j7FqSftn0R8ae55ZtUMleRRs53NnFCKmBtAfPYC3Y0EOQI6xfrOprKS3B2CZ15Y
I2TvFG4q0px9Gw0dZsqfHHQg9EMLEC2pBq+C/2QDGuVEtgfQ5/n5pLFC+aLUZ0A6
1KFCDE+CCsPUnCUw9oE5GztEnNttC07vmpqnT7U/xIX6yjeCb5xu55b02LmQ0eiv
pY54uAoIxi2uOQgBq7TknZcNjdMc7HJZpztjWzTw4nmdf9cn/MqA1oCGjWCvEwdF
MFmBhKB14buLYs9PF3/izy2T3w9o5r9Kxv5FPWis8cN6N6+MTELfdRdnMnixgBn5
uQKlt1FHydxGcKlUqzR+eo3yeVr3DSSeWdLQtdndS+RqNCOolJZOKyiyEzIRAdAk
BKHKPm4ubGoVJSY6+k1l5PRVfo2iz/AS9YMd5kbKxYfY+/c748FNcS7yVBdQSsFu
dreo3EdnGX5Fe0ox05guwutar+M+RVtfxABjnyTm5D8U/p5zh6kSblViXyh0sqaj
lPkJeeumLaN57l6v0oIHPKHTHRcWUuFz7oB9SEoTLkJWrpj1z4ayaTqYrKKRJS/C
/MUM0rWXqblu+q0lkp1KnsPXmh7AIIJJtF6vKe/tpb9gNh1biUje8ESr0v6h5T0A
SLKP9BeFPvkB3pv9GiURb3tsG2DHr/JARcaevBWtMYxbk1Dtnwc17F6OZSFm/bxY
g9vWLxiHc/YPfwQJZN1eQDLfZXGtSUe+q1WmfB17uWkmsaqC2mVa3hw8Plsc4fi5
HYgfzx78sCT9d4o75+2g8WjFhfuD07OBXsd24V1raG/6mubfpNpd1EWIFea0TEyC
BYDBCFrbx1hmQp2yAS54SqgIEWkEhJUL+gMjFw/MV45ASHtt14T31Ny/hgnPcKzK
YSv3+UZ4mY1yKUkNSDVVOIGGnyXyp1npLVsws/nowjbUtnQPgmQ8T3XgD4bXWvsr
0hDSBEZVqn8G52Z5se/PdO1xfeRa0f0qHbik6wwDntP7mNZB9SsT4Dvna3626AYa
iU26+X+dI23iLJISEss1iBt5uUig7L83PSw7TFO3C204ISEqfnk1MdCaGyfTQi5r
SznW9uhv1Eyd/dd5u+0wO/0b0CjY3ouvg9FEvps5T7IbA67ZgX3BFBReeY04gPNH
lwfRa/jIlXg93I7dvlLtqRvROVmCaI/OwylQCJyc+SxoUdfSVvMKT9y2l8q+Fdc9
MT0CaTB2bYp42yw8TpbyDFkayxbk3k5r8VAtEIDjyd9mAe1teJdHicRipsipzLhc
wcvXZ5US3uPcr2UuWwVxpBAzuRDGtWx9zcpLVQ4oRwSHQSA8FocZrKXWtRJmpSMu
BIT6mZRDnfoAXrfaJfqfpwynA+s1+smRV+/CXi5vJpo9pnBYX3vJvkA7I4g8Cc+l
5P0QC13wgNrTgOA6HBVGdSUDtIj4QjRoLy5q+swyVGVb0HjdaKiMMQCLa8Y20zGy
LAilFdCU+XUNeAYsGQDxQrC8TjcmEHmviIo1SVNaQ6UdNuK2unRe5JOls5ENHNqU
QhCct/c8T5Kgyjj0yVuLmVIwxQ3nHk1oMLZmZ2W6xt7uVSABPqRBnYp2y7I1687a
J/XSiEQsuA8ii1MZV5b3CL8vipMBGi1aCcTRU6dyheIAP0v/bufo5lEHgDy+fvEw
12Wr/OeK/+GvNLhGSLrLZ/N4y5McA3u1mnnLj2KYaXxB7tVQoLMAYMC/X0lnzLij
oiQTmC0L6TqZYYhigZvYNFZUy3R+8OvdMh//Y6Uo6fE+er2zBZDbUyrnmT+CfSDx
wkfeEAaseTmkXSJhqypewQaVDY9HFqTTeodEaBWXsRSUZflz15pIDN1FRgYOGCSW
h25DEpZctOftywxoOv/WG7L00Pa3nUP0uO7H6sJziTTbXqjAZ1DlTeId+ClRc/o/
l7gCqddnHYsMDdboMguEo8E0X1PqDieos3S5vcLFvqPsWP2vQU3s24jNVKrTWncl
85tHyFHh3tH8MZ7h2yFhT9UKFCq4wqBXL8rSYX0clfXZpXmMZdFJsziHICdzvB8X
q68mjrEeD9iQ4SuLgSI1GiQK8WZAy2SR2IAzoIx0jG6lT6sUp9rF7gkMPVNftqco
laQcbDGh8O/31XOrmFHMBk+JTA07DkvGD37pJl3HBEqRH8qGxSMsK6Sk2tN7NuZF
LZlaoDacSxncu2nl2uItFsdHo6U4XnfW9QfWxFjkHBRcJL/pbjmkWKBRkiG+bPx7
8kUkjTJqD8EYq7V4vc607XkvbtJSKNzfqYcsEqwA+DgrdXfjDynd2st5h1gFqS9J
5O3nscEG5cR3gj6ootwIcCCS6flPPNSJbrkJlua+9AytBH5eWYBR5agusHAq3DnU
jxmMP3aVKi0cCJSsCIbPXA7aaWJ7c3WEk579gMZk47NnLJkGEprz8/7ABsWT+mZ8
wAfzCrgTHkr6r96cGatdx1q3geoZsMnQQpkfq1Ign4A+417Nu5qhVm94b7eO5lVU
5RI1RhE4LClWpU2FLWymRr4Dw0HNohivQxXQuHsX3/sMOYLT3oU59eI8+dl7lRa8
WY7jmQoxAUOO0KQ8W0aQw4kGZy1BFzGlGb9uSoKTgV6bny4CDU3WwSFFu7Y1/Xn8
96hTXUYxFkc8gjtzdmJSY+g8eBFCUPICRfg9ax8A11rPQfqzB/RfHEsW9VbCzewM
Ania5V1xnlfldm1R412P++Z0XFnXSFPRZCKs2pV7glpnaXfiOsvMxwfTfzmQhSjw
Z82t8lRaDNQgxKTVx0PSZ3+CKbBB8tODokownCspoKi2cFWKa+rl38iwsZ2g6Eb3
y6eX9VMpqFrmKslmkYfIPT9uYdEadc/sF7tq8/ka+VaqopsDpszq5EYPaudUDLF9
7HLQj8KuX3tj5sqetiB3oCj9Dq8lQhnPJ8gJ295FAbxP3YCU3sgPzDxCndsNTUCP
rtGFu4OuxoWL94d+1PfOrxhGQ2KS0KZE4uZqO9KRk8y1nsep7PVD/T89gBWocLTR
6emfBlDuXoW9oOIjMu2/GtxquYVbbVJtOLjFowtLfXuB0iVS81YjSmVITmih25Om
vFxnHC3UoTwrQCTuHTn2fD2nSj4hBtmJi76NmUUkeChQ0O9XjYkl2yYZNj562+pF
p7ICOGM+/oExYw3wLdMRc50MRxJ7cQtWq+ph5SVVBSPjFBryqCGiofxn2qHKeGFZ
pfofV6Y8nGOwwmbPvMyV5HceCRGjHOOSY/yCbwmuXSEDDJvErxRqynFfEzxHH0Fk
ja1Ztev86cPDPeCSBsxMrxxXkWHhGgpjSASwDwFQH30BaTHESf7vii6+hNi7dJnP
EWjeipC0hKNjY1F2Yw7m9m0MLMrkyoattlWgjlT7ewaND0gB0mlfx6a04SjOvqWk
0NJvErkgG3XMr+0Hb8D4BIcgzS/6zdQTc49lCMC0G/dBLwslbI8shiDNDFjZMT+0
tuHqY+z8NB7Dz4Ezo9OCglp9dTENF5kjGasBkkyaFCW6yQ4kCzBnJ03tmSu5iUjN
729OX0WYcNvN0PxP4ip9GuzZfMIKED4DqAXf5dd/gZVwMksYmMuOmnsB/6EA/5tY
OX/PkJjaX6qGBzl7PeaL9YfvAKVcj4XeoE+Mr90+pVkaTdaGJ+wZiCzax0vxGA9g
x1GFMntzrBqtT4Q4Bpxk6TgQ9F0xtsOtwf91WE9mo+h+ttNdKcph/e3uo2XPJ+6Y
eP0ALBg2gGiBfev+5H1hNoYr9s1+EAOE6xyxgLcDUXm1gBJfx4SvUxE3KRrSaXx1
SbIZhSeU/pN3GFzvqR9iKwRH7Ed1rK0kpLm63L6IgDpXIiZ+9cTITaM1TtNpny96
lYRrysen9bCbwgyHagtNw7tuFS5Zhvyzw0RSp3g41DwWKKvmaLDa4ZdTeEez+nly
31ENW/Qt/OdZLTDpkQEs+i6G7JqWj9CEYVxqP/ZnO48kylYr0U/fHe0yHGWoy2yD
CtsBbrOKXssRIyEj6qYIw5jxQPNM7vT+rOsyZAra7Sil+PShWeeuNi/CxDxSk6gW
jxa+anh/qp3sTxAuONEho2yHYFF836pIs1dKUOx5QzT10s4/fdB1/Mjg8irGqhbw
qsHzbTDTOxbdaebWSPvAvnOYSwnlwB1bkVdrj4US4hg2TowaWpU/o8SUuh5HtDg3
FFpG5rn6lhNRuy7O1Q6eTa0ZOPvMDXhGzi8gZqmkbAq8U9bq6lETTo110f4ZynLO
Hydu+cvdh9zf55XGn8sjYggIItdLF4Rm/8nqelU7K+h39S5ilgedlFjvly4DJ6/k
o5Kv+Q1qJU38SaQ3M+dyWTXZ3cLER9B8PYmOxmpIqD2Dfh7KABDR/2S6MoKBKuA/
Fnjketc5gZpNmM+Ti0Ug0p380SEtrbpAnOl5E+5As/ty73IhJLhn5aBTfrv4+Ft+
qQ0E9oBfgc6GyiWSwHXyWX8JviKFRxdYauqkLpU94An3ITQ34BLABhcu/R9kA8JW
Zisf0nIId8DcejdlTAfPkfyvzVnG3DR19oeMQcYiSJ5fBd9iaQdID8e+HbqP4dHx
0OomseW2Amq3efR5rNdak0E6YNWCbAFBV+Vbx4sxtWbUIhYZjZDsPKl+Ox4k+4Zm
J8/+8CvW+EbMMz9wD39XpAWa+H8ygnHGr08zovrmU6H2d2q5x6EIDFFwhI/1fPzb
di32gjezFhiUFws/Kni5Nzv2Lfm9ybuoZ5DiQD++pbpNO7F1c3Vs5V0ShNWOzv3t
or7uR9DdAD+IoZybQX8azilra9A8gPDe4P1/QdYKaqasA1uky029E/+g0mBsw1Q5
ExRU+EHaAlartxDELQPJ07SuYD5EkbYmp7A2vqpTSGOT8mz6BQJ4DC2KGuV7fZYR
aUhw3B9JQ/seJRtrKso2UL4iXvOo8LILY1l5o27oXrpQUseZV9SC7A9g13PgmVC2
RGdYcRbImXSIWfnkKnio+lHufZd9xDkAAR39zc5PZufGDpnHj5UTWovh9b6vnTB7
rkKSRem4IxRsOCoUrmSDFRMLvn5beMiOolLtP+79eZbOBIQA3VDj+/8XiwVQ5tjx
vGiuW8NYbSeFuhjWj9EN+s5d0rE1vLfCe3Urdl/4N+8iaUKBF/jg320NJCB1Ggoe
c91tAD+HwwGMr8nnqy95RPVw0W8bcC5BuMG+YbftM+myv7xMiZAbbQvr3CzuYOhw
YfLGL9CUkUDQ8AiXM6Y33l0vaAIUW+d0FIW+ElsDxPNgH/a2/eBU1/addA5MDvP1
AHXrhKgQemROhyFFhl7XMNEhZZk3QKbBq+xTk8sSk2ytb22XPGH9fk+CuFnMv7NS
V5Kpb90LuAyz6OQkrFZPaEr7Rp9ftTo1vsXiBVldI/SlZAoVneYnYEk+YJO6z6CX
vrJNYYjpUCfaC+6wbVSdAdFiBDFiIkvIu3948OCl5sa8c9w87eXyHm/jxIYplvh2
9aQ1fulMiCfq5LdKdFDkvAuNYTwmqPowtqXW6irvZ2fysNcxYHUVUnhIjL7Njfhw
wWxjkr35xPg7exWhwq1dsxptNozc5EA43mSMAyoNMTPteNrhWpkn90aeLWlCwr/F
CvjQ60ezL3cM+ixanpYu5HDB53EBoJ+V6SCT6Xdi8QtL1sStHYhSzqEr/+lBwaeI
THNcPbyaXhXSZ2+2v9DS75donpofkoFvZiDDKXgo4o4gBXdtuom6LRufRK+2C0cg
7c/YQqkQ8efHAUlM3Qb/MJiKO11rz0RyBum+JNV9aEDK5kYFYfD6442csINiO7iC
xfH5AquE6CQdATfiNa4eoUHKKOtiC4JfrbCXYtOkv3qiyV9V7WRtC+tSt4elqZmh
PCJbN6Ooz7yArSb2umxSvS+Om9O7KQcr3BbDsUwNfLZZka+y0jUr7Opy2aEUKHo5
4RAiLKvlOtub/MtakDrz8gMl31lgOkBqLkPayu+0v5lTADZMjGpUvYcpSq2UPhIk
OK4jGSUSSJipLMWZaMpg8dFxD2D5nZVwodrPgOQYX5g589540OJ3sFT4v2YQVFPe
ax9mhWGquG0HFAE1bD3l84Lzc6OwuDymFqi5vzW53AqcDdZTXxFL0mzd7xdAnsJo
f1fekOun+WLmCCp+V2Y6n5jth1TGSzAWL5hlfOM74w8x0By/hxkvhIXcfk6k5w9Y
2/5EQedQZ9s8/fySBCKluTTljQ8zHf9kwNTvifVv3vLnoYT/8J0CA4RQY9OuJh6T
m/H8rezghaaQdzgztRjp+986Z2o3eDqR1AzGcybX2/FDWB/KK6SITBaVTbs6Aelf
NIVZ8KAcuZ4nJERLH9mIn/wXPXmHoypWaEWFdr67srn5vgfBBJiE7Yf84Nmof3wd
DHgDOEYLiBvB5WRqIn+XMwRVMi5Qt+cHDcxEcgbaGXGWqkPqwvp76MVNDlvD00vJ
NyGELyg9p2Bh7QTZIv53SIqnXovmUexEDsxAPnF5FN0xqIenDxCneS5IuKlHRJTB
`protect END_PROTECTED
