-- HostSystem.vhd

-- Generated using ACDS version 13.0sp1 232 at 2021.04.18.19:44:09

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity HostSystem is
	port (
		clk_clk       : in std_logic := '0'; --   clk.clk
		reset_reset_n : in std_logic := '0'  -- reset.reset_n
	);
end entity HostSystem;

architecture rtl of HostSystem is
	component HostSystem_memory is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(63 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X'              -- reset_req
		);
	end component HostSystem_memory;

	component HostSystem_cpu is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			d_address     : out std_logic_vector(13 downto 0);                    -- address
			d_byteenable  : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read        : out std_logic;                                        -- read
			d_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			d_write       : out std_logic;                                        -- write
			d_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			i_address     : out std_logic_vector(13 downto 0);                    -- address
			i_read        : out std_logic;                                        -- read
			i_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			d_irq         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			no_ci_readra  : out std_logic                                         -- readra
		);
	end component HostSystem_cpu;

	component reg32_avalon_interface is
		port (
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write_en   : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			add        : in  std_logic                     := 'X';             -- address
			read_en    : in  std_logic                     := 'X';             -- read
			chipselect : in  std_logic                     := 'X';             -- chipselect
			clock      : in  std_logic                     := 'X';             -- clk
			resetn     : in  std_logic                     := 'X'              -- reset_n
		);
	end component reg32_avalon_interface;

	component altera_merlin_master_agent is
		generic (
			PKT_PROTECTION_H          : integer := 80;
			PKT_PROTECTION_L          : integer := 80;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_BURSTWRAP_H           : integer := 79;
			PKT_BURSTWRAP_L           : integer := 77;
			PKT_BURST_SIZE_H          : integer := 86;
			PKT_BURST_SIZE_L          : integer := 84;
			PKT_BURST_TYPE_H          : integer := 94;
			PKT_BURST_TYPE_L          : integer := 93;
			PKT_BYTE_CNT_H            : integer := 76;
			PKT_BYTE_CNT_L            : integer := 74;
			PKT_ADDR_H                : integer := 73;
			PKT_ADDR_L                : integer := 42;
			PKT_TRANS_COMPRESSED_READ : integer := 41;
			PKT_TRANS_POSTED          : integer := 40;
			PKT_TRANS_WRITE           : integer := 39;
			PKT_TRANS_READ            : integer := 38;
			PKT_TRANS_LOCK            : integer := 82;
			PKT_TRANS_EXCLUSIVE       : integer := 83;
			PKT_DATA_H                : integer := 37;
			PKT_DATA_L                : integer := 6;
			PKT_BYTEEN_H              : integer := 5;
			PKT_BYTEEN_L              : integer := 2;
			PKT_SRC_ID_H              : integer := 1;
			PKT_SRC_ID_L              : integer := 1;
			PKT_DEST_ID_H             : integer := 0;
			PKT_DEST_ID_L             : integer := 0;
			PKT_THREAD_ID_H           : integer := 88;
			PKT_THREAD_ID_L           : integer := 87;
			PKT_CACHE_H               : integer := 92;
			PKT_CACHE_L               : integer := 89;
			PKT_DATA_SIDEBAND_H       : integer := 105;
			PKT_DATA_SIDEBAND_L       : integer := 98;
			PKT_QOS_H                 : integer := 109;
			PKT_QOS_L                 : integer := 106;
			PKT_ADDR_SIDEBAND_H       : integer := 97;
			PKT_ADDR_SIDEBAND_L       : integer := 93;
			PKT_RESPONSE_STATUS_H     : integer := 111;
			PKT_RESPONSE_STATUS_L     : integer := 110;
			ST_DATA_W                 : integer := 112;
			ST_CHANNEL_W              : integer := 1;
			AV_BURSTCOUNT_W           : integer := 3;
			SUPPRESS_0_BYTEEN_RSP     : integer := 1;
			ID                        : integer := 1;
			BURSTWRAP_VALUE           : integer := 4;
			CACHE_VALUE               : integer := 0;
			SECURE_ACCESS_BIT         : integer := 1;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			av_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_write                : in  std_logic                     := 'X';             -- write
			av_read                 : in  std_logic                     := 'X';             -- read
			av_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest          : out std_logic;                                        -- waitrequest
			av_readdatavalid        : out std_logic;                                        -- readdatavalid
			av_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			av_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_lock                 : in  std_logic                     := 'X';             -- lock
			cp_valid                : out std_logic;                                        -- valid
			cp_data                 : out std_logic_vector(83 downto 0);                    -- data
			cp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_endofpacket          : out std_logic;                                        -- endofpacket
			cp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : in  std_logic                     := 'X';             -- valid
			rp_data                 : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			rp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			rp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			rp_ready                : out std_logic;                                        -- ready
			av_response             : out std_logic_vector(1 downto 0);                     -- response
			av_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid   : out std_logic                                         -- writeresponsevalid
		);
	end component altera_merlin_master_agent;

	component HostSystem_addr_router is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(83 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component HostSystem_addr_router;

	component HostSystem_id_router is
		port (
			sink_ready         : out std_logic;                                         -- ready
			sink_valid         : in  std_logic                      := 'X';             -- valid
			sink_data          : in  std_logic_vector(119 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                      := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                      := 'X';             -- endofpacket
			clk                : in  std_logic                      := 'X';             -- clk
			reset              : in  std_logic                      := 'X';             -- reset
			src_ready          : in  std_logic                      := 'X';             -- ready
			src_valid          : out std_logic;                                         -- valid
			src_data           : out std_logic_vector(119 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                      -- channel
			src_startofpacket  : out std_logic;                                         -- startofpacket
			src_endofpacket    : out std_logic                                          -- endofpacket
		);
	end component HostSystem_id_router;

	component HostSystem_id_router_001 is
		port (
			sink_ready         : out std_logic;                                        -- ready
			sink_valid         : in  std_logic                     := 'X';             -- valid
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			src_ready          : in  std_logic                     := 'X';             -- ready
			src_valid          : out std_logic;                                        -- valid
			src_data           : out std_logic_vector(83 downto 0);                    -- data
			src_channel        : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket  : out std_logic;                                        -- startofpacket
			src_endofpacket    : out std_logic                                         -- endofpacket
		);
	end component HostSystem_id_router_001;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS        : integer := 6;
			OUTPUT_RESET_SYNC_EDGES : string  := "deassert";
			SYNC_DEPTH              : integer := 2;
			RESET_REQUEST_PRESENT   : integer := 0
		);
		port (
			reset_in0  : in  std_logic := 'X'; -- reset
			clk        : in  std_logic := 'X'; -- clk
			reset_out  : out std_logic;        -- reset
			reset_req  : out std_logic;        -- reset_req
			reset_in1  : in  std_logic := 'X'; -- reset
			reset_in2  : in  std_logic := 'X'; -- reset
			reset_in3  : in  std_logic := 'X'; -- reset
			reset_in4  : in  std_logic := 'X'; -- reset
			reset_in5  : in  std_logic := 'X'; -- reset
			reset_in6  : in  std_logic := 'X'; -- reset
			reset_in7  : in  std_logic := 'X'; -- reset
			reset_in8  : in  std_logic := 'X'; -- reset
			reset_in9  : in  std_logic := 'X'; -- reset
			reset_in10 : in  std_logic := 'X'; -- reset
			reset_in11 : in  std_logic := 'X'; -- reset
			reset_in12 : in  std_logic := 'X'; -- reset
			reset_in13 : in  std_logic := 'X'; -- reset
			reset_in14 : in  std_logic := 'X'; -- reset
			reset_in15 : in  std_logic := 'X'  -- reset
		);
	end component altera_reset_controller;

	component HostSystem_cmd_xbar_demux is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			sink_ready         : out std_logic;                                        -- ready
			sink_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink_valid         : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- valid
			src0_ready         : in  std_logic                     := 'X';             -- ready
			src0_valid         : out std_logic;                                        -- valid
			src0_data          : out std_logic_vector(83 downto 0);                    -- data
			src0_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src0_startofpacket : out std_logic;                                        -- startofpacket
			src0_endofpacket   : out std_logic;                                        -- endofpacket
			src1_ready         : in  std_logic                     := 'X';             -- ready
			src1_valid         : out std_logic;                                        -- valid
			src1_data          : out std_logic_vector(83 downto 0);                    -- data
			src1_channel       : out std_logic_vector(1 downto 0);                     -- channel
			src1_startofpacket : out std_logic;                                        -- startofpacket
			src1_endofpacket   : out std_logic                                         -- endofpacket
		);
	end component HostSystem_cmd_xbar_demux;

	component HostSystem_cmd_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(83 downto 0);                    -- data
			src_channel         : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component HostSystem_cmd_xbar_mux;

	component HostSystem_rsp_xbar_mux is
		port (
			clk                 : in  std_logic                     := 'X';             -- clk
			reset               : in  std_logic                     := 'X';             -- reset
			src_ready           : in  std_logic                     := 'X';             -- ready
			src_valid           : out std_logic;                                        -- valid
			src_data            : out std_logic_vector(83 downto 0);                    -- data
			src_channel         : out std_logic_vector(1 downto 0);                     -- channel
			src_startofpacket   : out std_logic;                                        -- startofpacket
			src_endofpacket     : out std_logic;                                        -- endofpacket
			sink0_ready         : out std_logic;                                        -- ready
			sink0_valid         : in  std_logic                     := 'X';             -- valid
			sink0_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink0_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink0_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink0_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			sink1_ready         : out std_logic;                                        -- ready
			sink1_valid         : in  std_logic                     := 'X';             -- valid
			sink1_channel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			sink1_data          : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			sink1_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			sink1_endofpacket   : in  std_logic                     := 'X'              -- endofpacket
		);
	end component HostSystem_rsp_xbar_mux;

	component HostSystem_irq_mapper is
		port (
			clk        : in  std_logic                     := 'X'; -- clk
			reset      : in  std_logic                     := 'X'; -- reset
			sender_irq : out std_logic_vector(31 downto 0)         -- irq
		);
	end component HostSystem_irq_mapper;

	component hostsystem_memory_s1_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(63 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(63 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(9 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_readdata              : in  std_logic_vector(63 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(63 downto 0);                    -- writedata
			av_byteenable            : out std_logic_vector(7 downto 0);                     -- byteenable
			av_chipselect            : out std_logic;                                        -- chipselect
			av_clken                 : out std_logic;                                        -- clken
			av_read                  : out std_logic;                                        -- read
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(7 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component hostsystem_memory_s1_translator;

	component hostsystem_exemplo_novo_0_avalon_slave_0_translator is
		generic (
			AV_ADDRESS_W                   : integer := 30;
			AV_DATA_W                      : integer := 32;
			UAV_DATA_W                     : integer := 32;
			AV_BURSTCOUNT_W                : integer := 4;
			AV_BYTEENABLE_W                : integer := 4;
			UAV_BYTEENABLE_W               : integer := 4;
			UAV_ADDRESS_W                  : integer := 32;
			UAV_BURSTCOUNT_W               : integer := 4;
			AV_READLATENCY                 : integer := 0;
			USE_READDATAVALID              : integer := 1;
			USE_WAITREQUEST                : integer := 1;
			USE_UAV_CLKEN                  : integer := 0;
			USE_READRESPONSE               : integer := 0;
			USE_WRITERESPONSE              : integer := 0;
			AV_SYMBOLS_PER_WORD            : integer := 4;
			AV_ADDRESS_SYMBOLS             : integer := 0;
			AV_BURSTCOUNT_SYMBOLS          : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR     : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR    : integer := 0;
			AV_REQUIRE_UNALIGNED_ADDRESSES : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0;
			AV_READ_WAIT_CYCLES            : integer := 0;
			AV_WRITE_WAIT_CYCLES           : integer := 0;
			AV_SETUP_WAIT_CYCLES           : integer := 0;
			AV_DATA_HOLD_CYCLES            : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			uav_burstcount           : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			uav_read                 : in  std_logic                     := 'X';             -- read
			uav_write                : in  std_logic                     := 'X';             -- write
			uav_waitrequest          : out std_logic;                                        -- waitrequest
			uav_readdatavalid        : out std_logic;                                        -- readdatavalid
			uav_byteenable           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			uav_readdata             : out std_logic_vector(31 downto 0);                    -- readdata
			uav_writedata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			uav_lock                 : in  std_logic                     := 'X';             -- lock
			uav_debugaccess          : in  std_logic                     := 'X';             -- debugaccess
			av_address               : out std_logic_vector(0 downto 0);                     -- address
			av_write                 : out std_logic;                                        -- write
			av_read                  : out std_logic;                                        -- read
			av_readdata              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			av_writedata             : out std_logic_vector(31 downto 0);                    -- writedata
			av_chipselect            : out std_logic;                                        -- chipselect
			av_begintransfer         : out std_logic;                                        -- begintransfer
			av_beginbursttransfer    : out std_logic;                                        -- beginbursttransfer
			av_burstcount            : out std_logic_vector(0 downto 0);                     -- burstcount
			av_byteenable            : out std_logic_vector(3 downto 0);                     -- byteenable
			av_readdatavalid         : in  std_logic                     := 'X';             -- readdatavalid
			av_waitrequest           : in  std_logic                     := 'X';             -- waitrequest
			av_writebyteenable       : out std_logic_vector(3 downto 0);                     -- writebyteenable
			av_lock                  : out std_logic;                                        -- lock
			av_clken                 : out std_logic;                                        -- clken
			uav_clken                : in  std_logic                     := 'X';             -- clken
			av_debugaccess           : out std_logic;                                        -- debugaccess
			av_outputenable          : out std_logic;                                        -- outputenable
			uav_response             : out std_logic_vector(1 downto 0);                     -- response
			av_response              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			uav_writeresponserequest : in  std_logic                     := 'X';             -- writeresponserequest
			uav_writeresponsevalid   : out std_logic;                                        -- writeresponsevalid
			av_writeresponserequest  : out std_logic;                                        -- writeresponserequest
			av_writeresponsevalid    : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component hostsystem_exemplo_novo_0_avalon_slave_0_translator;

	component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                      := 'X';             -- clk
			reset             : in  std_logic                      := 'X';             -- reset
			in_data           : in  std_logic_vector(120 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                      := 'X';             -- valid
			in_ready          : out std_logic;                                         -- ready
			in_startofpacket  : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                      := 'X';             -- endofpacket
			out_data          : out std_logic_vector(120 downto 0);                    -- data
			out_valid         : out std_logic;                                         -- valid
			out_ready         : in  std_logic                      := 'X';             -- ready
			out_startofpacket : out std_logic;                                         -- startofpacket
			out_endofpacket   : out std_logic;                                         -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- address
			csr_read          : in  std_logic                      := 'X';             -- read
			csr_write         : in  std_logic                      := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                     -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0)  := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                         -- data
			almost_empty_data : out std_logic;                                         -- data
			in_empty          : in  std_logic                      := 'X';             -- empty
			out_empty         : out std_logic;                                         -- empty
			in_error          : in  std_logic                      := 'X';             -- error
			out_error         : out std_logic;                                         -- error
			in_channel        : in  std_logic                      := 'X';             -- channel
			out_channel       : out std_logic                                          -- channel
		);
	end component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo is
		generic (
			SYMBOLS_PER_BEAT    : integer := 1;
			BITS_PER_SYMBOL     : integer := 8;
			FIFO_DEPTH          : integer := 16;
			CHANNEL_WIDTH       : integer := 0;
			ERROR_WIDTH         : integer := 0;
			USE_PACKETS         : integer := 0;
			USE_FILL_LEVEL      : integer := 0;
			EMPTY_LATENCY       : integer := 3;
			USE_MEMORY_BLOCKS   : integer := 1;
			USE_STORE_FORWARD   : integer := 0;
			USE_ALMOST_FULL_IF  : integer := 0;
			USE_ALMOST_EMPTY_IF : integer := 0
		);
		port (
			clk               : in  std_logic                     := 'X';             -- clk
			reset             : in  std_logic                     := 'X';             -- reset
			in_data           : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			in_valid          : in  std_logic                     := 'X';             -- valid
			in_ready          : out std_logic;                                        -- ready
			in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			out_data          : out std_logic_vector(84 downto 0);                    -- data
			out_valid         : out std_logic;                                        -- valid
			out_ready         : in  std_logic                     := 'X';             -- ready
			out_startofpacket : out std_logic;                                        -- startofpacket
			out_endofpacket   : out std_logic;                                        -- endofpacket
			csr_address       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			csr_read          : in  std_logic                     := 'X';             -- read
			csr_write         : in  std_logic                     := 'X';             -- write
			csr_readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			csr_writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			almost_full_data  : out std_logic;                                        -- data
			almost_empty_data : out std_logic;                                        -- data
			in_empty          : in  std_logic                     := 'X';             -- empty
			out_empty         : out std_logic;                                        -- empty
			in_error          : in  std_logic                     := 'X';             -- error
			out_error         : out std_logic;                                        -- error
			in_channel        : in  std_logic                     := 'X';             -- channel
			out_channel       : out std_logic                                         -- channel
		);
	end component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo;

	component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                      := 'X';             -- clk
			reset                   : in  std_logic                      := 'X';             -- reset
			m0_address              : out std_logic_vector(13 downto 0);                     -- address
			m0_burstcount           : out std_logic_vector(3 downto 0);                      -- burstcount
			m0_byteenable           : out std_logic_vector(7 downto 0);                      -- byteenable
			m0_debugaccess          : out std_logic;                                         -- debugaccess
			m0_lock                 : out std_logic;                                         -- lock
			m0_readdata             : in  std_logic_vector(63 downto 0)  := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                      := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                         -- read
			m0_waitrequest          : in  std_logic                      := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(63 downto 0);                     -- writedata
			m0_write                : out std_logic;                                         -- write
			rp_endofpacket          : out std_logic;                                         -- endofpacket
			rp_ready                : in  std_logic                      := 'X';             -- ready
			rp_valid                : out std_logic;                                         -- valid
			rp_data                 : out std_logic_vector(119 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                         -- startofpacket
			cp_ready                : out std_logic;                                         -- ready
			cp_valid                : in  std_logic                      := 'X';             -- valid
			cp_data                 : in  std_logic_vector(119 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                      := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                      := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                         -- ready
			rf_sink_valid           : in  std_logic                      := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                      := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                      := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(120 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                      := 'X';             -- ready
			rf_source_valid         : out std_logic;                                         -- valid
			rf_source_startofpacket : out std_logic;                                         -- startofpacket
			rf_source_endofpacket   : out std_logic;                                         -- endofpacket
			rf_source_data          : out std_logic_vector(120 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                         -- ready
			rdata_fifo_sink_valid   : in  std_logic                      := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(65 downto 0)  := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                      := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                         -- valid
			rdata_fifo_src_data     : out std_logic_vector(65 downto 0);                     -- data
			m0_response             : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                         -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                      := 'X'              -- writeresponsevalid
		);
	end component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent;

	component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent is
		generic (
			PKT_DATA_H                : integer := 31;
			PKT_DATA_L                : integer := 0;
			PKT_BEGIN_BURST           : integer := 81;
			PKT_SYMBOL_W              : integer := 8;
			PKT_BYTEEN_H              : integer := 71;
			PKT_BYTEEN_L              : integer := 68;
			PKT_ADDR_H                : integer := 63;
			PKT_ADDR_L                : integer := 32;
			PKT_TRANS_COMPRESSED_READ : integer := 67;
			PKT_TRANS_POSTED          : integer := 66;
			PKT_TRANS_WRITE           : integer := 65;
			PKT_TRANS_READ            : integer := 64;
			PKT_TRANS_LOCK            : integer := 87;
			PKT_SRC_ID_H              : integer := 74;
			PKT_SRC_ID_L              : integer := 72;
			PKT_DEST_ID_H             : integer := 77;
			PKT_DEST_ID_L             : integer := 75;
			PKT_BURSTWRAP_H           : integer := 85;
			PKT_BURSTWRAP_L           : integer := 82;
			PKT_BYTE_CNT_H            : integer := 81;
			PKT_BYTE_CNT_L            : integer := 78;
			PKT_PROTECTION_H          : integer := 86;
			PKT_PROTECTION_L          : integer := 86;
			PKT_RESPONSE_STATUS_H     : integer := 89;
			PKT_RESPONSE_STATUS_L     : integer := 88;
			PKT_BURST_SIZE_H          : integer := 92;
			PKT_BURST_SIZE_L          : integer := 90;
			ST_CHANNEL_W              : integer := 8;
			ST_DATA_W                 : integer := 93;
			AVS_BURSTCOUNT_W          : integer := 4;
			SUPPRESS_0_BYTEEN_CMD     : integer := 1;
			PREVENT_FIFO_OVERFLOW     : integer := 0;
			USE_READRESPONSE          : integer := 0;
			USE_WRITERESPONSE         : integer := 0
		);
		port (
			clk                     : in  std_logic                     := 'X';             -- clk
			reset                   : in  std_logic                     := 'X';             -- reset
			m0_address              : out std_logic_vector(13 downto 0);                    -- address
			m0_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			m0_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			m0_debugaccess          : out std_logic;                                        -- debugaccess
			m0_lock                 : out std_logic;                                        -- lock
			m0_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			m0_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			m0_read                 : out std_logic;                                        -- read
			m0_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			m0_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			m0_write                : out std_logic;                                        -- write
			rp_endofpacket          : out std_logic;                                        -- endofpacket
			rp_ready                : in  std_logic                     := 'X';             -- ready
			rp_valid                : out std_logic;                                        -- valid
			rp_data                 : out std_logic_vector(83 downto 0);                    -- data
			rp_startofpacket        : out std_logic;                                        -- startofpacket
			cp_ready                : out std_logic;                                        -- ready
			cp_valid                : in  std_logic                     := 'X';             -- valid
			cp_data                 : in  std_logic_vector(83 downto 0) := (others => 'X'); -- data
			cp_startofpacket        : in  std_logic                     := 'X';             -- startofpacket
			cp_endofpacket          : in  std_logic                     := 'X';             -- endofpacket
			cp_channel              : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- channel
			rf_sink_ready           : out std_logic;                                        -- ready
			rf_sink_valid           : in  std_logic                     := 'X';             -- valid
			rf_sink_startofpacket   : in  std_logic                     := 'X';             -- startofpacket
			rf_sink_endofpacket     : in  std_logic                     := 'X';             -- endofpacket
			rf_sink_data            : in  std_logic_vector(84 downto 0) := (others => 'X'); -- data
			rf_source_ready         : in  std_logic                     := 'X';             -- ready
			rf_source_valid         : out std_logic;                                        -- valid
			rf_source_startofpacket : out std_logic;                                        -- startofpacket
			rf_source_endofpacket   : out std_logic;                                        -- endofpacket
			rf_source_data          : out std_logic_vector(84 downto 0);                    -- data
			rdata_fifo_sink_ready   : out std_logic;                                        -- ready
			rdata_fifo_sink_valid   : in  std_logic                     := 'X';             -- valid
			rdata_fifo_sink_data    : in  std_logic_vector(33 downto 0) := (others => 'X'); -- data
			rdata_fifo_src_ready    : in  std_logic                     := 'X';             -- ready
			rdata_fifo_src_valid    : out std_logic;                                        -- valid
			rdata_fifo_src_data     : out std_logic_vector(33 downto 0);                    -- data
			m0_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			m0_writeresponserequest : out std_logic;                                        -- writeresponserequest
			m0_writeresponsevalid   : in  std_logic                     := 'X'              -- writeresponsevalid
		);
	end component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent;

	component hostsystem_width_adapter is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(83 downto 0)  := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(119 downto 0);                    -- data
			out_channel          : out std_logic_vector(1 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component hostsystem_width_adapter;

	component hostsystem_width_adapter_001 is
		generic (
			IN_PKT_ADDR_H                 : integer := 60;
			IN_PKT_ADDR_L                 : integer := 36;
			IN_PKT_DATA_H                 : integer := 31;
			IN_PKT_DATA_L                 : integer := 0;
			IN_PKT_BYTEEN_H               : integer := 35;
			IN_PKT_BYTEEN_L               : integer := 32;
			IN_PKT_BYTE_CNT_H             : integer := 63;
			IN_PKT_BYTE_CNT_L             : integer := 61;
			IN_PKT_TRANS_COMPRESSED_READ  : integer := 65;
			IN_PKT_BURSTWRAP_H            : integer := 67;
			IN_PKT_BURSTWRAP_L            : integer := 66;
			IN_PKT_BURST_SIZE_H           : integer := 70;
			IN_PKT_BURST_SIZE_L           : integer := 68;
			IN_PKT_RESPONSE_STATUS_H      : integer := 72;
			IN_PKT_RESPONSE_STATUS_L      : integer := 71;
			IN_PKT_TRANS_EXCLUSIVE        : integer := 73;
			IN_PKT_BURST_TYPE_H           : integer := 75;
			IN_PKT_BURST_TYPE_L           : integer := 74;
			IN_ST_DATA_W                  : integer := 76;
			OUT_PKT_ADDR_H                : integer := 60;
			OUT_PKT_ADDR_L                : integer := 36;
			OUT_PKT_DATA_H                : integer := 31;
			OUT_PKT_DATA_L                : integer := 0;
			OUT_PKT_BYTEEN_H              : integer := 35;
			OUT_PKT_BYTEEN_L              : integer := 32;
			OUT_PKT_BYTE_CNT_H            : integer := 63;
			OUT_PKT_BYTE_CNT_L            : integer := 61;
			OUT_PKT_TRANS_COMPRESSED_READ : integer := 65;
			OUT_PKT_BURST_SIZE_H          : integer := 68;
			OUT_PKT_BURST_SIZE_L          : integer := 66;
			OUT_PKT_RESPONSE_STATUS_H     : integer := 70;
			OUT_PKT_RESPONSE_STATUS_L     : integer := 69;
			OUT_PKT_TRANS_EXCLUSIVE       : integer := 71;
			OUT_PKT_BURST_TYPE_H          : integer := 73;
			OUT_PKT_BURST_TYPE_L          : integer := 72;
			OUT_ST_DATA_W                 : integer := 74;
			ST_CHANNEL_W                  : integer := 32;
			OPTIMIZE_FOR_RSP              : integer := 0;
			RESPONSE_PATH                 : integer := 0
		);
		port (
			clk                  : in  std_logic                      := 'X';             -- clk
			reset                : in  std_logic                      := 'X';             -- reset
			in_valid             : in  std_logic                      := 'X';             -- valid
			in_channel           : in  std_logic_vector(1 downto 0)   := (others => 'X'); -- channel
			in_startofpacket     : in  std_logic                      := 'X';             -- startofpacket
			in_endofpacket       : in  std_logic                      := 'X';             -- endofpacket
			in_ready             : out std_logic;                                         -- ready
			in_data              : in  std_logic_vector(119 downto 0) := (others => 'X'); -- data
			out_endofpacket      : out std_logic;                                         -- endofpacket
			out_data             : out std_logic_vector(83 downto 0);                     -- data
			out_channel          : out std_logic_vector(1 downto 0);                      -- channel
			out_valid            : out std_logic;                                         -- valid
			out_ready            : in  std_logic                      := 'X';             -- ready
			out_startofpacket    : out std_logic;                                         -- startofpacket
			in_command_size_data : in  std_logic_vector(2 downto 0)   := (others => 'X')  -- data
		);
	end component hostsystem_width_adapter_001;

	component hostsystem_cpu_instruction_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(13 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component hostsystem_cpu_instruction_master_translator;

	component hostsystem_cpu_data_master_translator is
		generic (
			AV_ADDRESS_W                : integer := 32;
			AV_DATA_W                   : integer := 32;
			AV_BURSTCOUNT_W             : integer := 4;
			AV_BYTEENABLE_W             : integer := 4;
			UAV_ADDRESS_W               : integer := 38;
			UAV_BURSTCOUNT_W            : integer := 10;
			USE_READ                    : integer := 1;
			USE_WRITE                   : integer := 1;
			USE_BEGINBURSTTRANSFER      : integer := 0;
			USE_BEGINTRANSFER           : integer := 0;
			USE_CHIPSELECT              : integer := 0;
			USE_BURSTCOUNT              : integer := 1;
			USE_READDATAVALID           : integer := 1;
			USE_WAITREQUEST             : integer := 1;
			USE_READRESPONSE            : integer := 0;
			USE_WRITERESPONSE           : integer := 0;
			AV_SYMBOLS_PER_WORD         : integer := 4;
			AV_ADDRESS_SYMBOLS          : integer := 0;
			AV_BURSTCOUNT_SYMBOLS       : integer := 0;
			AV_CONSTANT_BURST_BEHAVIOR  : integer := 0;
			UAV_CONSTANT_BURST_BEHAVIOR : integer := 0;
			AV_LINEWRAPBURSTS           : integer := 0;
			AV_REGISTERINCOMINGSIGNALS  : integer := 0
		);
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			uav_address              : out std_logic_vector(13 downto 0);                    -- address
			uav_burstcount           : out std_logic_vector(2 downto 0);                     -- burstcount
			uav_read                 : out std_logic;                                        -- read
			uav_write                : out std_logic;                                        -- write
			uav_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			uav_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			uav_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			uav_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			uav_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			uav_lock                 : out std_logic;                                        -- lock
			uav_debugaccess          : out std_logic;                                        -- debugaccess
			av_address               : in  std_logic_vector(13 downto 0) := (others => 'X'); -- address
			av_waitrequest           : out std_logic;                                        -- waitrequest
			av_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			av_read                  : in  std_logic                     := 'X';             -- read
			av_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			av_write                 : in  std_logic                     := 'X';             -- write
			av_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_burstcount            : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- burstcount
			av_beginbursttransfer    : in  std_logic                     := 'X';             -- beginbursttransfer
			av_begintransfer         : in  std_logic                     := 'X';             -- begintransfer
			av_chipselect            : in  std_logic                     := 'X';             -- chipselect
			av_readdatavalid         : out std_logic;                                        -- readdatavalid
			av_lock                  : in  std_logic                     := 'X';             -- lock
			av_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			uav_clken                : out std_logic;                                        -- clken
			av_clken                 : in  std_logic                     := 'X';             -- clken
			uav_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			av_response              : out std_logic_vector(1 downto 0);                     -- response
			uav_writeresponserequest : out std_logic;                                        -- writeresponserequest
			uav_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			av_writeresponserequest  : in  std_logic                     := 'X';             -- writeresponserequest
			av_writeresponsevalid    : out std_logic                                         -- writeresponsevalid
		);
	end component hostsystem_cpu_data_master_translator;

	signal cpu_instruction_master_waitrequest                                                                 : std_logic;                      -- cpu_instruction_master_translator:av_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                                                     : std_logic_vector(13 downto 0);  -- cpu:i_address -> cpu_instruction_master_translator:av_address
	signal cpu_instruction_master_read                                                                        : std_logic;                      -- cpu:i_read -> cpu_instruction_master_translator:av_read
	signal cpu_instruction_master_readdata                                                                    : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:av_readdata -> cpu:i_readdata
	signal cpu_data_master_waitrequest                                                                        : std_logic;                      -- cpu_data_master_translator:av_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_writedata                                                                          : std_logic_vector(31 downto 0);  -- cpu:d_writedata -> cpu_data_master_translator:av_writedata
	signal cpu_data_master_address                                                                            : std_logic_vector(13 downto 0);  -- cpu:d_address -> cpu_data_master_translator:av_address
	signal cpu_data_master_write                                                                              : std_logic;                      -- cpu:d_write -> cpu_data_master_translator:av_write
	signal cpu_data_master_read                                                                               : std_logic;                      -- cpu:d_read -> cpu_data_master_translator:av_read
	signal cpu_data_master_readdata                                                                           : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:av_readdata -> cpu:d_readdata
	signal cpu_data_master_byteenable                                                                         : std_logic_vector(3 downto 0);   -- cpu:d_byteenable -> cpu_data_master_translator:av_byteenable
	signal memory_s1_translator_avalon_anti_slave_0_writedata                                                 : std_logic_vector(63 downto 0);  -- memory_s1_translator:av_writedata -> memory:writedata
	signal memory_s1_translator_avalon_anti_slave_0_address                                                   : std_logic_vector(9 downto 0);   -- memory_s1_translator:av_address -> memory:address
	signal memory_s1_translator_avalon_anti_slave_0_chipselect                                                : std_logic;                      -- memory_s1_translator:av_chipselect -> memory:chipselect
	signal memory_s1_translator_avalon_anti_slave_0_clken                                                     : std_logic;                      -- memory_s1_translator:av_clken -> memory:clken
	signal memory_s1_translator_avalon_anti_slave_0_write                                                     : std_logic;                      -- memory_s1_translator:av_write -> memory:write
	signal memory_s1_translator_avalon_anti_slave_0_readdata                                                  : std_logic_vector(63 downto 0);  -- memory:readdata -> memory_s1_translator:av_readdata
	signal memory_s1_translator_avalon_anti_slave_0_byteenable                                                : std_logic_vector(7 downto 0);   -- memory_s1_translator:av_byteenable -> memory:byteenable
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata                             : std_logic_vector(31 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator:av_writedata -> exemplo_novo_0:writedata
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_address                               : std_logic_vector(0 downto 0);   -- exemplo_novo_0_avalon_slave_0_translator:av_address -> exemplo_novo_0:add
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect                            : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator:av_chipselect -> exemplo_novo_0:chipselect
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_write                                 : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator:av_write -> exemplo_novo_0:write_en
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_read                                  : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator:av_read -> exemplo_novo_0:read_en
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata                              : std_logic_vector(31 downto 0);  -- exemplo_novo_0:readdata -> exemplo_novo_0_avalon_slave_0_translator:av_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_waitrequest                            : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_instruction_master_translator:uav_waitrequest
	signal cpu_instruction_master_translator_avalon_universal_master_0_burstcount                             : std_logic_vector(2 downto 0);   -- cpu_instruction_master_translator:uav_burstcount -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_instruction_master_translator_avalon_universal_master_0_writedata                              : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator:uav_writedata -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_instruction_master_translator_avalon_universal_master_0_address                                : std_logic_vector(13 downto 0);  -- cpu_instruction_master_translator:uav_address -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_instruction_master_translator_avalon_universal_master_0_lock                                   : std_logic;                      -- cpu_instruction_master_translator:uav_lock -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_instruction_master_translator_avalon_universal_master_0_write                                  : std_logic;                      -- cpu_instruction_master_translator:uav_write -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_instruction_master_translator_avalon_universal_master_0_read                                   : std_logic;                      -- cpu_instruction_master_translator:uav_read -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdata                               : std_logic_vector(31 downto 0);  -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_instruction_master_translator:uav_readdata
	signal cpu_instruction_master_translator_avalon_universal_master_0_debugaccess                            : std_logic;                      -- cpu_instruction_master_translator:uav_debugaccess -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_instruction_master_translator_avalon_universal_master_0_byteenable                             : std_logic_vector(3 downto 0);   -- cpu_instruction_master_translator:uav_byteenable -> cpu_instruction_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid                          : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_instruction_master_translator:uav_readdatavalid
	signal cpu_data_master_translator_avalon_universal_master_0_waitrequest                                   : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_waitrequest -> cpu_data_master_translator:uav_waitrequest
	signal cpu_data_master_translator_avalon_universal_master_0_burstcount                                    : std_logic_vector(2 downto 0);   -- cpu_data_master_translator:uav_burstcount -> cpu_data_master_translator_avalon_universal_master_0_agent:av_burstcount
	signal cpu_data_master_translator_avalon_universal_master_0_writedata                                     : std_logic_vector(31 downto 0);  -- cpu_data_master_translator:uav_writedata -> cpu_data_master_translator_avalon_universal_master_0_agent:av_writedata
	signal cpu_data_master_translator_avalon_universal_master_0_address                                       : std_logic_vector(13 downto 0);  -- cpu_data_master_translator:uav_address -> cpu_data_master_translator_avalon_universal_master_0_agent:av_address
	signal cpu_data_master_translator_avalon_universal_master_0_lock                                          : std_logic;                      -- cpu_data_master_translator:uav_lock -> cpu_data_master_translator_avalon_universal_master_0_agent:av_lock
	signal cpu_data_master_translator_avalon_universal_master_0_write                                         : std_logic;                      -- cpu_data_master_translator:uav_write -> cpu_data_master_translator_avalon_universal_master_0_agent:av_write
	signal cpu_data_master_translator_avalon_universal_master_0_read                                          : std_logic;                      -- cpu_data_master_translator:uav_read -> cpu_data_master_translator_avalon_universal_master_0_agent:av_read
	signal cpu_data_master_translator_avalon_universal_master_0_readdata                                      : std_logic_vector(31 downto 0);  -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdata -> cpu_data_master_translator:uav_readdata
	signal cpu_data_master_translator_avalon_universal_master_0_debugaccess                                   : std_logic;                      -- cpu_data_master_translator:uav_debugaccess -> cpu_data_master_translator_avalon_universal_master_0_agent:av_debugaccess
	signal cpu_data_master_translator_avalon_universal_master_0_byteenable                                    : std_logic_vector(3 downto 0);   -- cpu_data_master_translator:uav_byteenable -> cpu_data_master_translator_avalon_universal_master_0_agent:av_byteenable
	signal cpu_data_master_translator_avalon_universal_master_0_readdatavalid                                 : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> cpu_data_master_translator:uav_readdatavalid
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest                                 : std_logic;                      -- memory_s1_translator:uav_waitrequest -> memory_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount                                  : std_logic_vector(3 downto 0);   -- memory_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> memory_s1_translator:uav_burstcount
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata                                   : std_logic_vector(63 downto 0);  -- memory_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> memory_s1_translator:uav_writedata
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_address                                     : std_logic_vector(13 downto 0);  -- memory_s1_translator_avalon_universal_slave_0_agent:m0_address -> memory_s1_translator:uav_address
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_write                                       : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:m0_write -> memory_s1_translator:uav_write
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_lock                                        : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:m0_lock -> memory_s1_translator:uav_lock
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_read                                        : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:m0_read -> memory_s1_translator:uav_read
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata                                    : std_logic_vector(63 downto 0);  -- memory_s1_translator:uav_readdata -> memory_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid                               : std_logic;                      -- memory_s1_translator:uav_readdatavalid -> memory_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess                                 : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> memory_s1_translator:uav_debugaccess
	signal memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable                                  : std_logic_vector(7 downto 0);   -- memory_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> memory_s1_translator:uav_byteenable
	signal memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket                          : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid                                : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket                        : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data                                 : std_logic_vector(120 downto 0); -- memory_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready                                : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> memory_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket                       : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid                             : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket                     : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data                              : std_logic_vector(120 downto 0); -- memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready                             : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid                           : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data                            : std_logic_vector(65 downto 0);  -- memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready                           : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> memory_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest             : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator:uav_waitrequest -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount              : std_logic_vector(2 downto 0);   -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> exemplo_novo_0_avalon_slave_0_translator:uav_burstcount
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata               : std_logic_vector(31 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> exemplo_novo_0_avalon_slave_0_translator:uav_writedata
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address                 : std_logic_vector(13 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> exemplo_novo_0_avalon_slave_0_translator:uav_address
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write                   : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> exemplo_novo_0_avalon_slave_0_translator:uav_write
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock                    : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> exemplo_novo_0_avalon_slave_0_translator:uav_lock
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read                    : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> exemplo_novo_0_avalon_slave_0_translator:uav_read
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata                : std_logic_vector(31 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator:uav_readdata -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid           : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator:uav_readdatavalid -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess             : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> exemplo_novo_0_avalon_slave_0_translator:uav_debugaccess
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable              : std_logic_vector(3 downto 0);   -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> exemplo_novo_0_avalon_slave_0_translator:uav_byteenable
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket      : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid            : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket    : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data             : std_logic_vector(84 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready            : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket   : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid         : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data          : std_logic_vector(84 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready         : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid       : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data        : std_logic_vector(33 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready       : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket                   : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid                         : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket                 : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data                          : std_logic_vector(83 downto 0);  -- cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	signal cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready                         : std_logic;                      -- addr_router:sink_ready -> cpu_instruction_master_translator_avalon_universal_master_0_agent:cp_ready
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket                          : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_001:sink_endofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid                                : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_001:sink_valid
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket                        : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_001:sink_startofpacket
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_data                                 : std_logic_vector(83 downto 0);  -- cpu_data_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_001:sink_data
	signal cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready                                : std_logic;                      -- addr_router_001:sink_ready -> cpu_data_master_translator_avalon_universal_master_0_agent:cp_ready
	signal memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket                                 : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rp_valid                                       : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	signal memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket                               : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	signal memory_s1_translator_avalon_universal_slave_0_agent_rp_data                                        : std_logic_vector(119 downto 0); -- memory_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	signal memory_s1_translator_avalon_universal_slave_0_agent_rp_ready                                       : std_logic;                      -- id_router:sink_ready -> memory_s1_translator_avalon_universal_slave_0_agent:rp_ready
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket             : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid                   : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket           : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data                    : std_logic_vector(83 downto 0);  -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	signal exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready                   : std_logic;                      -- id_router_001:sink_ready -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	signal rst_controller_reset_out_reset                                                                     : std_logic;                      -- rst_controller:reset_out -> [addr_router:reset, addr_router_001:reset, cmd_xbar_demux:reset, cmd_xbar_demux_001:reset, cmd_xbar_mux:reset, cmd_xbar_mux_001:reset, cpu_data_master_translator:reset, cpu_data_master_translator_avalon_universal_master_0_agent:reset, cpu_instruction_master_translator:reset, cpu_instruction_master_translator_avalon_universal_master_0_agent:reset, exemplo_novo_0_avalon_slave_0_translator:reset, exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, irq_mapper:reset, memory:reset, memory_s1_translator:reset, memory_s1_translator_avalon_universal_slave_0_agent:reset, memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux:reset, rsp_xbar_mux_001:reset, rst_controller_reset_out_reset:in, width_adapter:reset, width_adapter_001:reset]
	signal rst_controller_reset_out_reset_req                                                                 : std_logic;                      -- rst_controller:reset_req -> memory:reset_req
	signal cmd_xbar_demux_src0_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux:src0_endofpacket -> cmd_xbar_mux:sink0_endofpacket
	signal cmd_xbar_demux_src0_valid                                                                          : std_logic;                      -- cmd_xbar_demux:src0_valid -> cmd_xbar_mux:sink0_valid
	signal cmd_xbar_demux_src0_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux:src0_startofpacket -> cmd_xbar_mux:sink0_startofpacket
	signal cmd_xbar_demux_src0_data                                                                           : std_logic_vector(83 downto 0);  -- cmd_xbar_demux:src0_data -> cmd_xbar_mux:sink0_data
	signal cmd_xbar_demux_src0_channel                                                                        : std_logic_vector(1 downto 0);   -- cmd_xbar_demux:src0_channel -> cmd_xbar_mux:sink0_channel
	signal cmd_xbar_demux_src0_ready                                                                          : std_logic;                      -- cmd_xbar_mux:sink0_ready -> cmd_xbar_demux:src0_ready
	signal cmd_xbar_demux_src1_endofpacket                                                                    : std_logic;                      -- cmd_xbar_demux:src1_endofpacket -> cmd_xbar_mux_001:sink0_endofpacket
	signal cmd_xbar_demux_src1_valid                                                                          : std_logic;                      -- cmd_xbar_demux:src1_valid -> cmd_xbar_mux_001:sink0_valid
	signal cmd_xbar_demux_src1_startofpacket                                                                  : std_logic;                      -- cmd_xbar_demux:src1_startofpacket -> cmd_xbar_mux_001:sink0_startofpacket
	signal cmd_xbar_demux_src1_data                                                                           : std_logic_vector(83 downto 0);  -- cmd_xbar_demux:src1_data -> cmd_xbar_mux_001:sink0_data
	signal cmd_xbar_demux_src1_channel                                                                        : std_logic_vector(1 downto 0);   -- cmd_xbar_demux:src1_channel -> cmd_xbar_mux_001:sink0_channel
	signal cmd_xbar_demux_src1_ready                                                                          : std_logic;                      -- cmd_xbar_mux_001:sink0_ready -> cmd_xbar_demux:src1_ready
	signal cmd_xbar_demux_001_src0_endofpacket                                                                : std_logic;                      -- cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux:sink1_endofpacket
	signal cmd_xbar_demux_001_src0_valid                                                                      : std_logic;                      -- cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux:sink1_valid
	signal cmd_xbar_demux_001_src0_startofpacket                                                              : std_logic;                      -- cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux:sink1_startofpacket
	signal cmd_xbar_demux_001_src0_data                                                                       : std_logic_vector(83 downto 0);  -- cmd_xbar_demux_001:src0_data -> cmd_xbar_mux:sink1_data
	signal cmd_xbar_demux_001_src0_channel                                                                    : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux:sink1_channel
	signal cmd_xbar_demux_001_src0_ready                                                                      : std_logic;                      -- cmd_xbar_mux:sink1_ready -> cmd_xbar_demux_001:src0_ready
	signal cmd_xbar_demux_001_src1_endofpacket                                                                : std_logic;                      -- cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_001:sink1_endofpacket
	signal cmd_xbar_demux_001_src1_valid                                                                      : std_logic;                      -- cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_001:sink1_valid
	signal cmd_xbar_demux_001_src1_startofpacket                                                              : std_logic;                      -- cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_001:sink1_startofpacket
	signal cmd_xbar_demux_001_src1_data                                                                       : std_logic_vector(83 downto 0);  -- cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_001:sink1_data
	signal cmd_xbar_demux_001_src1_channel                                                                    : std_logic_vector(1 downto 0);   -- cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_001:sink1_channel
	signal cmd_xbar_demux_001_src1_ready                                                                      : std_logic;                      -- cmd_xbar_mux_001:sink1_ready -> cmd_xbar_demux_001:src1_ready
	signal rsp_xbar_demux_src0_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	signal rsp_xbar_demux_src0_valid                                                                          : std_logic;                      -- rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	signal rsp_xbar_demux_src0_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	signal rsp_xbar_demux_src0_data                                                                           : std_logic_vector(83 downto 0);  -- rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	signal rsp_xbar_demux_src0_channel                                                                        : std_logic_vector(1 downto 0);   -- rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	signal rsp_xbar_demux_src0_ready                                                                          : std_logic;                      -- rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	signal rsp_xbar_demux_src1_endofpacket                                                                    : std_logic;                      -- rsp_xbar_demux:src1_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	signal rsp_xbar_demux_src1_valid                                                                          : std_logic;                      -- rsp_xbar_demux:src1_valid -> rsp_xbar_mux_001:sink0_valid
	signal rsp_xbar_demux_src1_startofpacket                                                                  : std_logic;                      -- rsp_xbar_demux:src1_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	signal rsp_xbar_demux_src1_data                                                                           : std_logic_vector(83 downto 0);  -- rsp_xbar_demux:src1_data -> rsp_xbar_mux_001:sink0_data
	signal rsp_xbar_demux_src1_channel                                                                        : std_logic_vector(1 downto 0);   -- rsp_xbar_demux:src1_channel -> rsp_xbar_mux_001:sink0_channel
	signal rsp_xbar_demux_src1_ready                                                                          : std_logic;                      -- rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux:src1_ready
	signal rsp_xbar_demux_001_src0_endofpacket                                                                : std_logic;                      -- rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	signal rsp_xbar_demux_001_src0_valid                                                                      : std_logic;                      -- rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	signal rsp_xbar_demux_001_src0_startofpacket                                                              : std_logic;                      -- rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	signal rsp_xbar_demux_001_src0_data                                                                       : std_logic_vector(83 downto 0);  -- rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	signal rsp_xbar_demux_001_src0_channel                                                                    : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	signal rsp_xbar_demux_001_src0_ready                                                                      : std_logic;                      -- rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	signal rsp_xbar_demux_001_src1_endofpacket                                                                : std_logic;                      -- rsp_xbar_demux_001:src1_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	signal rsp_xbar_demux_001_src1_valid                                                                      : std_logic;                      -- rsp_xbar_demux_001:src1_valid -> rsp_xbar_mux_001:sink1_valid
	signal rsp_xbar_demux_001_src1_startofpacket                                                              : std_logic;                      -- rsp_xbar_demux_001:src1_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	signal rsp_xbar_demux_001_src1_data                                                                       : std_logic_vector(83 downto 0);  -- rsp_xbar_demux_001:src1_data -> rsp_xbar_mux_001:sink1_data
	signal rsp_xbar_demux_001_src1_channel                                                                    : std_logic_vector(1 downto 0);   -- rsp_xbar_demux_001:src1_channel -> rsp_xbar_mux_001:sink1_channel
	signal rsp_xbar_demux_001_src1_ready                                                                      : std_logic;                      -- rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_001:src1_ready
	signal addr_router_src_endofpacket                                                                        : std_logic;                      -- addr_router:src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	signal addr_router_src_valid                                                                              : std_logic;                      -- addr_router:src_valid -> cmd_xbar_demux:sink_valid
	signal addr_router_src_startofpacket                                                                      : std_logic;                      -- addr_router:src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	signal addr_router_src_data                                                                               : std_logic_vector(83 downto 0);  -- addr_router:src_data -> cmd_xbar_demux:sink_data
	signal addr_router_src_channel                                                                            : std_logic_vector(1 downto 0);   -- addr_router:src_channel -> cmd_xbar_demux:sink_channel
	signal addr_router_src_ready                                                                              : std_logic;                      -- cmd_xbar_demux:sink_ready -> addr_router:src_ready
	signal rsp_xbar_mux_src_endofpacket                                                                       : std_logic;                      -- rsp_xbar_mux:src_endofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_src_valid                                                                             : std_logic;                      -- rsp_xbar_mux:src_valid -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_src_startofpacket                                                                     : std_logic;                      -- rsp_xbar_mux:src_startofpacket -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_src_data                                                                              : std_logic_vector(83 downto 0);  -- rsp_xbar_mux:src_data -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_src_channel                                                                           : std_logic_vector(1 downto 0);   -- rsp_xbar_mux:src_channel -> cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_src_ready                                                                             : std_logic;                      -- cpu_instruction_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux:src_ready
	signal addr_router_001_src_endofpacket                                                                    : std_logic;                      -- addr_router_001:src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	signal addr_router_001_src_valid                                                                          : std_logic;                      -- addr_router_001:src_valid -> cmd_xbar_demux_001:sink_valid
	signal addr_router_001_src_startofpacket                                                                  : std_logic;                      -- addr_router_001:src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	signal addr_router_001_src_data                                                                           : std_logic_vector(83 downto 0);  -- addr_router_001:src_data -> cmd_xbar_demux_001:sink_data
	signal addr_router_001_src_channel                                                                        : std_logic_vector(1 downto 0);   -- addr_router_001:src_channel -> cmd_xbar_demux_001:sink_channel
	signal addr_router_001_src_ready                                                                          : std_logic;                      -- cmd_xbar_demux_001:sink_ready -> addr_router_001:src_ready
	signal rsp_xbar_mux_001_src_endofpacket                                                                   : std_logic;                      -- rsp_xbar_mux_001:src_endofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	signal rsp_xbar_mux_001_src_valid                                                                         : std_logic;                      -- rsp_xbar_mux_001:src_valid -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_valid
	signal rsp_xbar_mux_001_src_startofpacket                                                                 : std_logic;                      -- rsp_xbar_mux_001:src_startofpacket -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	signal rsp_xbar_mux_001_src_data                                                                          : std_logic_vector(83 downto 0);  -- rsp_xbar_mux_001:src_data -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_data
	signal rsp_xbar_mux_001_src_channel                                                                       : std_logic_vector(1 downto 0);   -- rsp_xbar_mux_001:src_channel -> cpu_data_master_translator_avalon_universal_master_0_agent:rp_channel
	signal rsp_xbar_mux_001_src_ready                                                                         : std_logic;                      -- cpu_data_master_translator_avalon_universal_master_0_agent:rp_ready -> rsp_xbar_mux_001:src_ready
	signal cmd_xbar_mux_001_src_endofpacket                                                                   : std_logic;                      -- cmd_xbar_mux_001:src_endofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal cmd_xbar_mux_001_src_valid                                                                         : std_logic;                      -- cmd_xbar_mux_001:src_valid -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	signal cmd_xbar_mux_001_src_startofpacket                                                                 : std_logic;                      -- cmd_xbar_mux_001:src_startofpacket -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal cmd_xbar_mux_001_src_data                                                                          : std_logic_vector(83 downto 0);  -- cmd_xbar_mux_001:src_data -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	signal cmd_xbar_mux_001_src_channel                                                                       : std_logic_vector(1 downto 0);   -- cmd_xbar_mux_001:src_channel -> exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	signal cmd_xbar_mux_001_src_ready                                                                         : std_logic;                      -- exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_mux_001:src_ready
	signal id_router_001_src_endofpacket                                                                      : std_logic;                      -- id_router_001:src_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	signal id_router_001_src_valid                                                                            : std_logic;                      -- id_router_001:src_valid -> rsp_xbar_demux_001:sink_valid
	signal id_router_001_src_startofpacket                                                                    : std_logic;                      -- id_router_001:src_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	signal id_router_001_src_data                                                                             : std_logic_vector(83 downto 0);  -- id_router_001:src_data -> rsp_xbar_demux_001:sink_data
	signal id_router_001_src_channel                                                                          : std_logic_vector(1 downto 0);   -- id_router_001:src_channel -> rsp_xbar_demux_001:sink_channel
	signal id_router_001_src_ready                                                                            : std_logic;                      -- rsp_xbar_demux_001:sink_ready -> id_router_001:src_ready
	signal cmd_xbar_mux_src_endofpacket                                                                       : std_logic;                      -- cmd_xbar_mux:src_endofpacket -> width_adapter:in_endofpacket
	signal cmd_xbar_mux_src_valid                                                                             : std_logic;                      -- cmd_xbar_mux:src_valid -> width_adapter:in_valid
	signal cmd_xbar_mux_src_startofpacket                                                                     : std_logic;                      -- cmd_xbar_mux:src_startofpacket -> width_adapter:in_startofpacket
	signal cmd_xbar_mux_src_data                                                                              : std_logic_vector(83 downto 0);  -- cmd_xbar_mux:src_data -> width_adapter:in_data
	signal cmd_xbar_mux_src_channel                                                                           : std_logic_vector(1 downto 0);   -- cmd_xbar_mux:src_channel -> width_adapter:in_channel
	signal cmd_xbar_mux_src_ready                                                                             : std_logic;                      -- width_adapter:in_ready -> cmd_xbar_mux:src_ready
	signal width_adapter_src_endofpacket                                                                      : std_logic;                      -- width_adapter:out_endofpacket -> memory_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	signal width_adapter_src_valid                                                                            : std_logic;                      -- width_adapter:out_valid -> memory_s1_translator_avalon_universal_slave_0_agent:cp_valid
	signal width_adapter_src_startofpacket                                                                    : std_logic;                      -- width_adapter:out_startofpacket -> memory_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	signal width_adapter_src_data                                                                             : std_logic_vector(119 downto 0); -- width_adapter:out_data -> memory_s1_translator_avalon_universal_slave_0_agent:cp_data
	signal width_adapter_src_ready                                                                            : std_logic;                      -- memory_s1_translator_avalon_universal_slave_0_agent:cp_ready -> width_adapter:out_ready
	signal width_adapter_src_channel                                                                          : std_logic_vector(1 downto 0);   -- width_adapter:out_channel -> memory_s1_translator_avalon_universal_slave_0_agent:cp_channel
	signal id_router_src_endofpacket                                                                          : std_logic;                      -- id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	signal id_router_src_valid                                                                                : std_logic;                      -- id_router:src_valid -> width_adapter_001:in_valid
	signal id_router_src_startofpacket                                                                        : std_logic;                      -- id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	signal id_router_src_data                                                                                 : std_logic_vector(119 downto 0); -- id_router:src_data -> width_adapter_001:in_data
	signal id_router_src_channel                                                                              : std_logic_vector(1 downto 0);   -- id_router:src_channel -> width_adapter_001:in_channel
	signal id_router_src_ready                                                                                : std_logic;                      -- width_adapter_001:in_ready -> id_router:src_ready
	signal width_adapter_001_src_endofpacket                                                                  : std_logic;                      -- width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	signal width_adapter_001_src_valid                                                                        : std_logic;                      -- width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	signal width_adapter_001_src_startofpacket                                                                : std_logic;                      -- width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	signal width_adapter_001_src_data                                                                         : std_logic_vector(83 downto 0);  -- width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	signal width_adapter_001_src_ready                                                                        : std_logic;                      -- rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	signal width_adapter_001_src_channel                                                                      : std_logic_vector(1 downto 0);   -- width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	signal cpu_d_irq_irq                                                                                      : std_logic_vector(31 downto 0);  -- irq_mapper:sender_irq -> cpu:d_irq
	signal reset_reset_n_ports_inv                                                                            : std_logic;                      -- reset_reset_n:inv -> rst_controller:reset_in0
	signal rst_controller_reset_out_reset_ports_inv                                                           : std_logic;                      -- rst_controller_reset_out_reset:inv -> [cpu:reset_n, exemplo_novo_0:resetn]

begin

	memory : component HostSystem_memory
		port map (
			clk        => clk_clk,                                             --   clk1.clk
			address    => memory_s1_translator_avalon_anti_slave_0_address,    --     s1.address
			clken      => memory_s1_translator_avalon_anti_slave_0_clken,      --       .clken
			chipselect => memory_s1_translator_avalon_anti_slave_0_chipselect, --       .chipselect
			write      => memory_s1_translator_avalon_anti_slave_0_write,      --       .write
			readdata   => memory_s1_translator_avalon_anti_slave_0_readdata,   --       .readdata
			writedata  => memory_s1_translator_avalon_anti_slave_0_writedata,  --       .writedata
			byteenable => memory_s1_translator_avalon_anti_slave_0_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,                      -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req                   --       .reset_req
		);

	cpu : component HostSystem_cpu
		port map (
			clk           => clk_clk,                                  --                       clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv, --                   reset_n.reset_n
			d_address     => cpu_data_master_address,                  --               data_master.address
			d_byteenable  => cpu_data_master_byteenable,               --                          .byteenable
			d_read        => cpu_data_master_read,                     --                          .read
			d_readdata    => cpu_data_master_readdata,                 --                          .readdata
			d_waitrequest => cpu_data_master_waitrequest,              --                          .waitrequest
			d_write       => cpu_data_master_write,                    --                          .write
			d_writedata   => cpu_data_master_writedata,                --                          .writedata
			i_address     => cpu_instruction_master_address,           --        instruction_master.address
			i_read        => cpu_instruction_master_read,              --                          .read
			i_readdata    => cpu_instruction_master_readdata,          --                          .readdata
			i_waitrequest => cpu_instruction_master_waitrequest,       --                          .waitrequest
			d_irq         => cpu_d_irq_irq,                            --                     d_irq.irq
			no_ci_readra  => open                                      -- custom_instruction_master.readra
		);

	exemplo_novo_0 : component reg32_avalon_interface
		port map (
			writedata  => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,  -- avalon_slave_0.writedata
			write_en   => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_write,      --               .write
			readdata   => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,   --               .readdata
			add        => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_address(0), --               .address
			read_en    => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_read,       --               .read
			chipselect => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect, --               .chipselect
			clock      => clk_clk,                                                                 --     clock_sink.clk
			resetn     => rst_controller_reset_out_reset_ports_inv                                 --     reset_sink.reset_n
		);

	cpu_instruction_master_translator : component hostsystem_cpu_instruction_master_translator
		generic map (
			AV_ADDRESS_W                => 14,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 14,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 0,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 1,
			AV_REGISTERINCOMINGSIGNALS  => 0
		)
		port map (
			clk                      => clk_clk,                                                                   --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                            --                     reset.reset
			uav_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_instruction_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_instruction_master_waitrequest,                                        --                          .waitrequest
			av_read                  => cpu_instruction_master_read,                                               --                          .read
			av_readdata              => cpu_instruction_master_readdata,                                           --                          .readdata
			av_burstcount            => "1",                                                                       --               (terminated)
			av_byteenable            => "1111",                                                                    --               (terminated)
			av_beginbursttransfer    => '0',                                                                       --               (terminated)
			av_begintransfer         => '0',                                                                       --               (terminated)
			av_chipselect            => '0',                                                                       --               (terminated)
			av_readdatavalid         => open,                                                                      --               (terminated)
			av_write                 => '0',                                                                       --               (terminated)
			av_writedata             => "00000000000000000000000000000000",                                        --               (terminated)
			av_lock                  => '0',                                                                       --               (terminated)
			av_debugaccess           => '0',                                                                       --               (terminated)
			uav_clken                => open,                                                                      --               (terminated)
			av_clken                 => '1',                                                                       --               (terminated)
			uav_response             => "00",                                                                      --               (terminated)
			av_response              => open,                                                                      --               (terminated)
			uav_writeresponserequest => open,                                                                      --               (terminated)
			uav_writeresponsevalid   => '0',                                                                       --               (terminated)
			av_writeresponserequest  => '0',                                                                       --               (terminated)
			av_writeresponsevalid    => open                                                                       --               (terminated)
		);

	cpu_data_master_translator : component hostsystem_cpu_data_master_translator
		generic map (
			AV_ADDRESS_W                => 14,
			AV_DATA_W                   => 32,
			AV_BURSTCOUNT_W             => 1,
			AV_BYTEENABLE_W             => 4,
			UAV_ADDRESS_W               => 14,
			UAV_BURSTCOUNT_W            => 3,
			USE_READ                    => 1,
			USE_WRITE                   => 1,
			USE_BEGINBURSTTRANSFER      => 0,
			USE_BEGINTRANSFER           => 0,
			USE_CHIPSELECT              => 0,
			USE_BURSTCOUNT              => 0,
			USE_READDATAVALID           => 0,
			USE_WAITREQUEST             => 1,
			USE_READRESPONSE            => 0,
			USE_WRITERESPONSE           => 0,
			AV_SYMBOLS_PER_WORD         => 4,
			AV_ADDRESS_SYMBOLS          => 1,
			AV_BURSTCOUNT_SYMBOLS       => 0,
			AV_CONSTANT_BURST_BEHAVIOR  => 0,
			UAV_CONSTANT_BURST_BEHAVIOR => 0,
			AV_LINEWRAPBURSTS           => 0,
			AV_REGISTERINCOMINGSIGNALS  => 1
		)
		port map (
			clk                      => clk_clk,                                                            --                       clk.clk
			reset                    => rst_controller_reset_out_reset,                                     --                     reset.reset
			uav_address              => cpu_data_master_translator_avalon_universal_master_0_address,       -- avalon_universal_master_0.address
			uav_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,    --                          .burstcount
			uav_read                 => cpu_data_master_translator_avalon_universal_master_0_read,          --                          .read
			uav_write                => cpu_data_master_translator_avalon_universal_master_0_write,         --                          .write
			uav_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,   --                          .waitrequest
			uav_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid, --                          .readdatavalid
			uav_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,    --                          .byteenable
			uav_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,      --                          .readdata
			uav_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,     --                          .writedata
			uav_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,          --                          .lock
			uav_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,   --                          .debugaccess
			av_address               => cpu_data_master_address,                                            --      avalon_anti_master_0.address
			av_waitrequest           => cpu_data_master_waitrequest,                                        --                          .waitrequest
			av_byteenable            => cpu_data_master_byteenable,                                         --                          .byteenable
			av_read                  => cpu_data_master_read,                                               --                          .read
			av_readdata              => cpu_data_master_readdata,                                           --                          .readdata
			av_write                 => cpu_data_master_write,                                              --                          .write
			av_writedata             => cpu_data_master_writedata,                                          --                          .writedata
			av_burstcount            => "1",                                                                --               (terminated)
			av_beginbursttransfer    => '0',                                                                --               (terminated)
			av_begintransfer         => '0',                                                                --               (terminated)
			av_chipselect            => '0',                                                                --               (terminated)
			av_readdatavalid         => open,                                                               --               (terminated)
			av_lock                  => '0',                                                                --               (terminated)
			av_debugaccess           => '0',                                                                --               (terminated)
			uav_clken                => open,                                                               --               (terminated)
			av_clken                 => '1',                                                                --               (terminated)
			uav_response             => "00",                                                               --               (terminated)
			av_response              => open,                                                               --               (terminated)
			uav_writeresponserequest => open,                                                               --               (terminated)
			uav_writeresponsevalid   => '0',                                                                --               (terminated)
			av_writeresponserequest  => '0',                                                                --               (terminated)
			av_writeresponsevalid    => open                                                                --               (terminated)
		);

	memory_s1_translator : component hostsystem_memory_s1_translator
		generic map (
			AV_ADDRESS_W                   => 10,
			AV_DATA_W                      => 64,
			UAV_DATA_W                     => 64,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 8,
			UAV_BYTEENABLE_W               => 8,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 4,
			AV_READLATENCY                 => 1,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 8,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 0,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                              --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                       --                    reset.reset
			uav_address              => memory_s1_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => memory_s1_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => memory_s1_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => memory_s1_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => memory_s1_translator_avalon_anti_slave_0_write,                       --                         .write
			av_readdata              => memory_s1_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => memory_s1_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_byteenable            => memory_s1_translator_avalon_anti_slave_0_byteenable,                  --                         .byteenable
			av_chipselect            => memory_s1_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_clken                 => memory_s1_translator_avalon_anti_slave_0_clken,                       --                         .clken
			av_read                  => open,                                                                 --              (terminated)
			av_begintransfer         => open,                                                                 --              (terminated)
			av_beginbursttransfer    => open,                                                                 --              (terminated)
			av_burstcount            => open,                                                                 --              (terminated)
			av_readdatavalid         => '0',                                                                  --              (terminated)
			av_waitrequest           => '0',                                                                  --              (terminated)
			av_writebyteenable       => open,                                                                 --              (terminated)
			av_lock                  => open,                                                                 --              (terminated)
			uav_clken                => '0',                                                                  --              (terminated)
			av_debugaccess           => open,                                                                 --              (terminated)
			av_outputenable          => open,                                                                 --              (terminated)
			uav_response             => open,                                                                 --              (terminated)
			av_response              => "00",                                                                 --              (terminated)
			uav_writeresponserequest => '0',                                                                  --              (terminated)
			uav_writeresponsevalid   => open,                                                                 --              (terminated)
			av_writeresponserequest  => open,                                                                 --              (terminated)
			av_writeresponsevalid    => '0'                                                                   --              (terminated)
		);

	exemplo_novo_0_avalon_slave_0_translator : component hostsystem_exemplo_novo_0_avalon_slave_0_translator
		generic map (
			AV_ADDRESS_W                   => 1,
			AV_DATA_W                      => 32,
			UAV_DATA_W                     => 32,
			AV_BURSTCOUNT_W                => 1,
			AV_BYTEENABLE_W                => 4,
			UAV_BYTEENABLE_W               => 4,
			UAV_ADDRESS_W                  => 14,
			UAV_BURSTCOUNT_W               => 3,
			AV_READLATENCY                 => 0,
			USE_READDATAVALID              => 0,
			USE_WAITREQUEST                => 0,
			USE_UAV_CLKEN                  => 0,
			USE_READRESPONSE               => 0,
			USE_WRITERESPONSE              => 0,
			AV_SYMBOLS_PER_WORD            => 4,
			AV_ADDRESS_SYMBOLS             => 0,
			AV_BURSTCOUNT_SYMBOLS          => 0,
			AV_CONSTANT_BURST_BEHAVIOR     => 0,
			UAV_CONSTANT_BURST_BEHAVIOR    => 0,
			AV_REQUIRE_UNALIGNED_ADDRESSES => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0,
			AV_READ_WAIT_CYCLES            => 1,
			AV_WRITE_WAIT_CYCLES           => 0,
			AV_SETUP_WAIT_CYCLES           => 0,
			AV_DATA_HOLD_CYCLES            => 0
		)
		port map (
			clk                      => clk_clk,                                                                                  --                      clk.clk
			reset                    => rst_controller_reset_out_reset,                                                           --                    reset.reset
			uav_address              => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,       -- avalon_universal_slave_0.address
			uav_burstcount           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,    --                         .burstcount
			uav_read                 => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,          --                         .read
			uav_write                => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,         --                         .write
			uav_waitrequest          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,   --                         .waitrequest
			uav_readdatavalid        => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid, --                         .readdatavalid
			uav_byteenable           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,    --                         .byteenable
			uav_readdata             => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,      --                         .readdata
			uav_writedata            => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,     --                         .writedata
			uav_lock                 => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,          --                         .lock
			uav_debugaccess          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,   --                         .debugaccess
			av_address               => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_address,                     --      avalon_anti_slave_0.address
			av_write                 => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_write,                       --                         .write
			av_read                  => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_read,                        --                         .read
			av_readdata              => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata,                    --                         .readdata
			av_writedata             => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata,                   --                         .writedata
			av_chipselect            => exemplo_novo_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect,                  --                         .chipselect
			av_begintransfer         => open,                                                                                     --              (terminated)
			av_beginbursttransfer    => open,                                                                                     --              (terminated)
			av_burstcount            => open,                                                                                     --              (terminated)
			av_byteenable            => open,                                                                                     --              (terminated)
			av_readdatavalid         => '0',                                                                                      --              (terminated)
			av_waitrequest           => '0',                                                                                      --              (terminated)
			av_writebyteenable       => open,                                                                                     --              (terminated)
			av_lock                  => open,                                                                                     --              (terminated)
			av_clken                 => open,                                                                                     --              (terminated)
			uav_clken                => '0',                                                                                      --              (terminated)
			av_debugaccess           => open,                                                                                     --              (terminated)
			av_outputenable          => open,                                                                                     --              (terminated)
			uav_response             => open,                                                                                     --              (terminated)
			av_response              => "00",                                                                                     --              (terminated)
			uav_writeresponserequest => '0',                                                                                      --              (terminated)
			uav_writeresponsevalid   => open,                                                                                     --              (terminated)
			av_writeresponserequest  => open,                                                                                     --              (terminated)
			av_writeresponsevalid    => '0'                                                                                       --              (terminated)
		);

	cpu_instruction_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_BEGIN_BURST           => 70,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			PKT_BURST_TYPE_H          => 67,
			PKT_BURST_TYPE_L          => 66,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 73,
			PKT_THREAD_ID_H           => 74,
			PKT_THREAD_ID_L           => 74,
			PKT_CACHE_H               => 81,
			PKT_CACHE_L               => 78,
			PKT_DATA_SIDEBAND_H       => 69,
			PKT_DATA_SIDEBAND_L       => 69,
			PKT_QOS_H                 => 71,
			PKT_QOS_L                 => 71,
			PKT_ADDR_SIDEBAND_H       => 68,
			PKT_ADDR_SIDEBAND_L       => 68,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			ST_DATA_W                 => 84,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 1,
			BURSTWRAP_VALUE           => 3,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                            --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			av_address              => cpu_instruction_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_instruction_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_instruction_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_instruction_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_instruction_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_instruction_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_instruction_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_instruction_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_instruction_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_instruction_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_instruction_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_src_valid,                                                             --        rp.valid
			rp_data                 => rsp_xbar_mux_src_data,                                                              --          .data
			rp_channel              => rsp_xbar_mux_src_channel,                                                           --          .channel
			rp_startofpacket        => rsp_xbar_mux_src_startofpacket,                                                     --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_src_endofpacket,                                                       --          .endofpacket
			rp_ready                => rsp_xbar_mux_src_ready,                                                             --          .ready
			av_response             => open,                                                                               -- (terminated)
			av_writeresponserequest => '0',                                                                                -- (terminated)
			av_writeresponsevalid   => open                                                                                -- (terminated)
		);

	cpu_data_master_translator_avalon_universal_master_0_agent : component altera_merlin_master_agent
		generic map (
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_BEGIN_BURST           => 70,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			PKT_BURST_TYPE_H          => 67,
			PKT_BURST_TYPE_L          => 66,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 56,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_TRANS_EXCLUSIVE       => 55,
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 73,
			PKT_THREAD_ID_H           => 74,
			PKT_THREAD_ID_L           => 74,
			PKT_CACHE_H               => 81,
			PKT_CACHE_L               => 78,
			PKT_DATA_SIDEBAND_H       => 69,
			PKT_DATA_SIDEBAND_L       => 69,
			PKT_QOS_H                 => 71,
			PKT_QOS_L                 => 71,
			PKT_ADDR_SIDEBAND_H       => 68,
			PKT_ADDR_SIDEBAND_L       => 68,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			ST_DATA_W                 => 84,
			ST_CHANNEL_W              => 2,
			AV_BURSTCOUNT_W           => 3,
			SUPPRESS_0_BYTEEN_RSP     => 1,
			ID                        => 0,
			BURSTWRAP_VALUE           => 7,
			CACHE_VALUE               => 0,
			SECURE_ACCESS_BIT         => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                     --       clk.clk
			reset                   => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			av_address              => cpu_data_master_translator_avalon_universal_master_0_address,                --        av.address
			av_write                => cpu_data_master_translator_avalon_universal_master_0_write,                  --          .write
			av_read                 => cpu_data_master_translator_avalon_universal_master_0_read,                   --          .read
			av_writedata            => cpu_data_master_translator_avalon_universal_master_0_writedata,              --          .writedata
			av_readdata             => cpu_data_master_translator_avalon_universal_master_0_readdata,               --          .readdata
			av_waitrequest          => cpu_data_master_translator_avalon_universal_master_0_waitrequest,            --          .waitrequest
			av_readdatavalid        => cpu_data_master_translator_avalon_universal_master_0_readdatavalid,          --          .readdatavalid
			av_byteenable           => cpu_data_master_translator_avalon_universal_master_0_byteenable,             --          .byteenable
			av_burstcount           => cpu_data_master_translator_avalon_universal_master_0_burstcount,             --          .burstcount
			av_debugaccess          => cpu_data_master_translator_avalon_universal_master_0_debugaccess,            --          .debugaccess
			av_lock                 => cpu_data_master_translator_avalon_universal_master_0_lock,                   --          .lock
			cp_valid                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --        cp.valid
			cp_data                 => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			cp_startofpacket        => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			cp_endofpacket          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			cp_ready                => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --          .ready
			rp_valid                => rsp_xbar_mux_001_src_valid,                                                  --        rp.valid
			rp_data                 => rsp_xbar_mux_001_src_data,                                                   --          .data
			rp_channel              => rsp_xbar_mux_001_src_channel,                                                --          .channel
			rp_startofpacket        => rsp_xbar_mux_001_src_startofpacket,                                          --          .startofpacket
			rp_endofpacket          => rsp_xbar_mux_001_src_endofpacket,                                            --          .endofpacket
			rp_ready                => rsp_xbar_mux_001_src_ready,                                                  --          .ready
			av_response             => open,                                                                        -- (terminated)
			av_writeresponserequest => '0',                                                                         -- (terminated)
			av_writeresponsevalid   => open                                                                         -- (terminated)
		);

	memory_s1_translator_avalon_universal_slave_0_agent : component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 63,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 106,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 71,
			PKT_BYTEEN_L              => 64,
			PKT_ADDR_H                => 85,
			PKT_ADDR_L                => 72,
			PKT_TRANS_COMPRESSED_READ => 86,
			PKT_TRANS_POSTED          => 87,
			PKT_TRANS_WRITE           => 88,
			PKT_TRANS_READ            => 89,
			PKT_TRANS_LOCK            => 90,
			PKT_SRC_ID_H              => 108,
			PKT_SRC_ID_L              => 108,
			PKT_DEST_ID_H             => 109,
			PKT_DEST_ID_L             => 109,
			PKT_BURSTWRAP_H           => 98,
			PKT_BURSTWRAP_L           => 96,
			PKT_BYTE_CNT_H            => 95,
			PKT_BYTE_CNT_L            => 92,
			PKT_PROTECTION_H          => 113,
			PKT_PROTECTION_L          => 111,
			PKT_RESPONSE_STATUS_H     => 119,
			PKT_RESPONSE_STATUS_L     => 118,
			PKT_BURST_SIZE_H          => 101,
			PKT_BURST_SIZE_L          => 99,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 120,
			AVS_BURSTCOUNT_W          => 4,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                        --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                 --       clk_reset.reset
			m0_address              => memory_s1_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => memory_s1_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => memory_s1_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => memory_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => memory_s1_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => memory_s1_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => memory_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => memory_s1_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => memory_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => memory_s1_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => memory_s1_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => memory_s1_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => width_adapter_src_ready,                                                        --              cp.ready
			cp_valid                => width_adapter_src_valid,                                                        --                .valid
			cp_data                 => width_adapter_src_data,                                                         --                .data
			cp_startofpacket        => width_adapter_src_startofpacket,                                                --                .startofpacket
			cp_endofpacket          => width_adapter_src_endofpacket,                                                  --                .endofpacket
			cp_channel              => width_adapter_src_channel,                                                      --                .channel
			rf_sink_ready           => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => memory_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                           --     (terminated)
			m0_writeresponserequest => open,                                                                           --     (terminated)
			m0_writeresponsevalid   => '0'                                                                             --     (terminated)
		);

	memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo : component hostsystem_memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 121,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                        --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                 -- clk_reset.reset
			in_data           => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => memory_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => memory_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                           -- (terminated)
			csr_read          => '0',                                                                            -- (terminated)
			csr_write         => '0',                                                                            -- (terminated)
			csr_readdata      => open,                                                                           -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                             -- (terminated)
			almost_full_data  => open,                                                                           -- (terminated)
			almost_empty_data => open,                                                                           -- (terminated)
			in_empty          => '0',                                                                            -- (terminated)
			out_empty         => open,                                                                           -- (terminated)
			in_error          => '0',                                                                            -- (terminated)
			out_error         => open,                                                                           -- (terminated)
			in_channel        => '0',                                                                            -- (terminated)
			out_channel       => open                                                                            -- (terminated)
		);

	exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent : component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent
		generic map (
			PKT_DATA_H                => 31,
			PKT_DATA_L                => 0,
			PKT_BEGIN_BURST           => 70,
			PKT_SYMBOL_W              => 8,
			PKT_BYTEEN_H              => 35,
			PKT_BYTEEN_L              => 32,
			PKT_ADDR_H                => 49,
			PKT_ADDR_L                => 36,
			PKT_TRANS_COMPRESSED_READ => 50,
			PKT_TRANS_POSTED          => 51,
			PKT_TRANS_WRITE           => 52,
			PKT_TRANS_READ            => 53,
			PKT_TRANS_LOCK            => 54,
			PKT_SRC_ID_H              => 72,
			PKT_SRC_ID_L              => 72,
			PKT_DEST_ID_H             => 73,
			PKT_DEST_ID_L             => 73,
			PKT_BURSTWRAP_H           => 62,
			PKT_BURSTWRAP_L           => 60,
			PKT_BYTE_CNT_H            => 59,
			PKT_BYTE_CNT_L            => 56,
			PKT_PROTECTION_H          => 77,
			PKT_PROTECTION_L          => 75,
			PKT_RESPONSE_STATUS_H     => 83,
			PKT_RESPONSE_STATUS_L     => 82,
			PKT_BURST_SIZE_H          => 65,
			PKT_BURST_SIZE_L          => 63,
			ST_CHANNEL_W              => 2,
			ST_DATA_W                 => 84,
			AVS_BURSTCOUNT_W          => 3,
			SUPPRESS_0_BYTEEN_CMD     => 0,
			PREVENT_FIFO_OVERFLOW     => 1,
			USE_READRESPONSE          => 0,
			USE_WRITERESPONSE         => 0
		)
		port map (
			clk                     => clk_clk,                                                                                            --             clk.clk
			reset                   => rst_controller_reset_out_reset,                                                                     --       clk_reset.reset
			m0_address              => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address,                 --              m0.address
			m0_burstcount           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount,              --                .burstcount
			m0_byteenable           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable,              --                .byteenable
			m0_debugaccess          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess,             --                .debugaccess
			m0_lock                 => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock,                    --                .lock
			m0_readdata             => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata,                --                .readdata
			m0_readdatavalid        => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid,           --                .readdatavalid
			m0_read                 => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read,                    --                .read
			m0_waitrequest          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest,             --                .waitrequest
			m0_writedata            => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata,               --                .writedata
			m0_write                => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write,                   --                .write
			rp_endofpacket          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,             --              rp.endofpacket
			rp_ready                => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,                   --                .ready
			rp_valid                => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,                   --                .valid
			rp_data                 => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,                    --                .data
			rp_startofpacket        => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket,           --                .startofpacket
			cp_ready                => cmd_xbar_mux_001_src_ready,                                                                         --              cp.ready
			cp_valid                => cmd_xbar_mux_001_src_valid,                                                                         --                .valid
			cp_data                 => cmd_xbar_mux_001_src_data,                                                                          --                .data
			cp_startofpacket        => cmd_xbar_mux_001_src_startofpacket,                                                                 --                .startofpacket
			cp_endofpacket          => cmd_xbar_mux_001_src_endofpacket,                                                                   --                .endofpacket
			cp_channel              => cmd_xbar_mux_001_src_channel,                                                                       --                .channel
			rf_sink_ready           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --         rf_sink.ready
			rf_sink_valid           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --                .valid
			rf_sink_startofpacket   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --                .startofpacket
			rf_sink_endofpacket     => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --                .endofpacket
			rf_sink_data            => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --                .data
			rf_source_ready         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --       rf_source.ready
			rf_source_valid         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --                .valid
			rf_source_startofpacket => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --                .startofpacket
			rf_source_endofpacket   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --                .endofpacket
			rf_source_data          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --                .data
			rdata_fifo_sink_ready   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       -- rdata_fifo_sink.ready
			rdata_fifo_sink_valid   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_sink_data    => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			rdata_fifo_src_ready    => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready,       --  rdata_fifo_src.ready
			rdata_fifo_src_valid    => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid,       --                .valid
			rdata_fifo_src_data     => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data,        --                .data
			m0_response             => "00",                                                                                               --     (terminated)
			m0_writeresponserequest => open,                                                                                               --     (terminated)
			m0_writeresponsevalid   => '0'                                                                                                 --     (terminated)
		);

	exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo : component hostsystem_exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo
		generic map (
			SYMBOLS_PER_BEAT    => 1,
			BITS_PER_SYMBOL     => 85,
			FIFO_DEPTH          => 2,
			CHANNEL_WIDTH       => 0,
			ERROR_WIDTH         => 0,
			USE_PACKETS         => 1,
			USE_FILL_LEVEL      => 0,
			EMPTY_LATENCY       => 1,
			USE_MEMORY_BLOCKS   => 0,
			USE_STORE_FORWARD   => 0,
			USE_ALMOST_FULL_IF  => 0,
			USE_ALMOST_EMPTY_IF => 0
		)
		port map (
			clk               => clk_clk,                                                                                            --       clk.clk
			reset             => rst_controller_reset_out_reset,                                                                     -- clk_reset.reset
			in_data           => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data,             --        in.data
			in_valid          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid,            --          .valid
			in_ready          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready,            --          .ready
			in_startofpacket  => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket,    --          .startofpacket
			in_endofpacket    => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket,      --          .endofpacket
			out_data          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data,          --       out.data
			out_valid         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid,         --          .valid
			out_ready         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready,         --          .ready
			out_startofpacket => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket, --          .startofpacket
			out_endofpacket   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket,   --          .endofpacket
			csr_address       => "00",                                                                                               -- (terminated)
			csr_read          => '0',                                                                                                -- (terminated)
			csr_write         => '0',                                                                                                -- (terminated)
			csr_readdata      => open,                                                                                               -- (terminated)
			csr_writedata     => "00000000000000000000000000000000",                                                                 -- (terminated)
			almost_full_data  => open,                                                                                               -- (terminated)
			almost_empty_data => open,                                                                                               -- (terminated)
			in_empty          => '0',                                                                                                -- (terminated)
			out_empty         => open,                                                                                               -- (terminated)
			in_error          => '0',                                                                                                -- (terminated)
			out_error         => open,                                                                                               -- (terminated)
			in_channel        => '0',                                                                                                -- (terminated)
			out_channel       => open                                                                                                -- (terminated)
		);

	addr_router : component HostSystem_addr_router
		port map (
			sink_ready         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_instruction_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                            --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                     -- clk_reset.reset
			src_ready          => addr_router_src_ready,                                                              --       src.ready
			src_valid          => addr_router_src_valid,                                                              --          .valid
			src_data           => addr_router_src_data,                                                               --          .data
			src_channel        => addr_router_src_channel,                                                            --          .channel
			src_startofpacket  => addr_router_src_startofpacket,                                                      --          .startofpacket
			src_endofpacket    => addr_router_src_endofpacket                                                         --          .endofpacket
		);

	addr_router_001 : component HostSystem_addr_router
		port map (
			sink_ready         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_ready,         --      sink.ready
			sink_valid         => cpu_data_master_translator_avalon_universal_master_0_agent_cp_valid,         --          .valid
			sink_data          => cpu_data_master_translator_avalon_universal_master_0_agent_cp_data,          --          .data
			sink_startofpacket => cpu_data_master_translator_avalon_universal_master_0_agent_cp_startofpacket, --          .startofpacket
			sink_endofpacket   => cpu_data_master_translator_avalon_universal_master_0_agent_cp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                     --       clk.clk
			reset              => rst_controller_reset_out_reset,                                              -- clk_reset.reset
			src_ready          => addr_router_001_src_ready,                                                   --       src.ready
			src_valid          => addr_router_001_src_valid,                                                   --          .valid
			src_data           => addr_router_001_src_data,                                                    --          .data
			src_channel        => addr_router_001_src_channel,                                                 --          .channel
			src_startofpacket  => addr_router_001_src_startofpacket,                                           --          .startofpacket
			src_endofpacket    => addr_router_001_src_endofpacket                                              --          .endofpacket
		);

	id_router : component HostSystem_id_router
		port map (
			sink_ready         => memory_s1_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => memory_s1_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => memory_s1_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => memory_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => memory_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                              --       clk.clk
			reset              => rst_controller_reset_out_reset,                                       -- clk_reset.reset
			src_ready          => id_router_src_ready,                                                  --       src.ready
			src_valid          => id_router_src_valid,                                                  --          .valid
			src_data           => id_router_src_data,                                                   --          .data
			src_channel        => id_router_src_channel,                                                --          .channel
			src_startofpacket  => id_router_src_startofpacket,                                          --          .startofpacket
			src_endofpacket    => id_router_src_endofpacket                                             --          .endofpacket
		);

	id_router_001 : component HostSystem_id_router_001
		port map (
			sink_ready         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready,         --      sink.ready
			sink_valid         => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid,         --          .valid
			sink_data          => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data,          --          .data
			sink_startofpacket => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket, --          .startofpacket
			sink_endofpacket   => exemplo_novo_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket,   --          .endofpacket
			clk                => clk_clk,                                                                                  --       clk.clk
			reset              => rst_controller_reset_out_reset,                                                           -- clk_reset.reset
			src_ready          => id_router_001_src_ready,                                                                  --       src.ready
			src_valid          => id_router_001_src_valid,                                                                  --          .valid
			src_data           => id_router_001_src_data,                                                                   --          .data
			src_channel        => id_router_001_src_channel,                                                                --          .channel
			src_startofpacket  => id_router_001_src_startofpacket,                                                          --          .startofpacket
			src_endofpacket    => id_router_001_src_endofpacket                                                             --          .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS        => 1,
			OUTPUT_RESET_SYNC_EDGES => "deassert",
			SYNC_DEPTH              => 2,
			RESET_REQUEST_PRESENT   => 1
		)
		port map (
			reset_in0  => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk        => clk_clk,                            --       clk.clk
			reset_out  => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req  => rst_controller_reset_out_reset_req, --          .reset_req
			reset_in1  => '0',                                -- (terminated)
			reset_in2  => '0',                                -- (terminated)
			reset_in3  => '0',                                -- (terminated)
			reset_in4  => '0',                                -- (terminated)
			reset_in5  => '0',                                -- (terminated)
			reset_in6  => '0',                                -- (terminated)
			reset_in7  => '0',                                -- (terminated)
			reset_in8  => '0',                                -- (terminated)
			reset_in9  => '0',                                -- (terminated)
			reset_in10 => '0',                                -- (terminated)
			reset_in11 => '0',                                -- (terminated)
			reset_in12 => '0',                                -- (terminated)
			reset_in13 => '0',                                -- (terminated)
			reset_in14 => '0',                                -- (terminated)
			reset_in15 => '0'                                 -- (terminated)
		);

	cmd_xbar_demux : component HostSystem_cmd_xbar_demux
		port map (
			clk                => clk_clk,                           --       clk.clk
			reset              => rst_controller_reset_out_reset,    -- clk_reset.reset
			sink_ready         => addr_router_src_ready,             --      sink.ready
			sink_channel       => addr_router_src_channel,           --          .channel
			sink_data          => addr_router_src_data,              --          .data
			sink_startofpacket => addr_router_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_demux_001 : component HostSystem_cmd_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => addr_router_001_src_ready,             --      sink.ready
			sink_channel       => addr_router_001_src_channel,           --          .channel
			sink_data          => addr_router_001_src_data,              --          .data
			sink_startofpacket => addr_router_001_src_startofpacket,     --          .startofpacket
			sink_endofpacket   => addr_router_001_src_endofpacket,       --          .endofpacket
			sink_valid(0)      => addr_router_001_src_valid,             --          .valid
			src0_ready         => cmd_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => cmd_xbar_demux_001_src0_data,          --          .data
			src0_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => cmd_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => cmd_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			src1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux : component HostSystem_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_src_ready,                --       src.ready
			src_valid           => cmd_xbar_mux_src_valid,                --          .valid
			src_data            => cmd_xbar_mux_src_data,                 --          .data
			src_channel         => cmd_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => cmd_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src0_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	cmd_xbar_mux_001 : component HostSystem_cmd_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => cmd_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => cmd_xbar_mux_001_src_valid,            --          .valid
			src_data            => cmd_xbar_mux_001_src_data,             --          .data
			src_channel         => cmd_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => cmd_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => cmd_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => cmd_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => cmd_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => cmd_xbar_demux_src1_channel,           --          .channel
			sink0_data          => cmd_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => cmd_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => cmd_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => cmd_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => cmd_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => cmd_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => cmd_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => cmd_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => cmd_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_demux : component HostSystem_cmd_xbar_demux
		port map (
			clk                => clk_clk,                             --       clk.clk
			reset              => rst_controller_reset_out_reset,      -- clk_reset.reset
			sink_ready         => width_adapter_001_src_ready,         --      sink.ready
			sink_channel       => width_adapter_001_src_channel,       --          .channel
			sink_data          => width_adapter_001_src_data,          --          .data
			sink_startofpacket => width_adapter_001_src_startofpacket, --          .startofpacket
			sink_endofpacket   => width_adapter_001_src_endofpacket,   --          .endofpacket
			sink_valid(0)      => width_adapter_001_src_valid,         --          .valid
			src0_ready         => rsp_xbar_demux_src0_ready,           --      src0.ready
			src0_valid         => rsp_xbar_demux_src0_valid,           --          .valid
			src0_data          => rsp_xbar_demux_src0_data,            --          .data
			src0_channel       => rsp_xbar_demux_src0_channel,         --          .channel
			src0_startofpacket => rsp_xbar_demux_src0_startofpacket,   --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_src0_endofpacket,     --          .endofpacket
			src1_ready         => rsp_xbar_demux_src1_ready,           --      src1.ready
			src1_valid         => rsp_xbar_demux_src1_valid,           --          .valid
			src1_data          => rsp_xbar_demux_src1_data,            --          .data
			src1_channel       => rsp_xbar_demux_src1_channel,         --          .channel
			src1_startofpacket => rsp_xbar_demux_src1_startofpacket,   --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_src1_endofpacket      --          .endofpacket
		);

	rsp_xbar_demux_001 : component HostSystem_cmd_xbar_demux
		port map (
			clk                => clk_clk,                               --       clk.clk
			reset              => rst_controller_reset_out_reset,        -- clk_reset.reset
			sink_ready         => id_router_001_src_ready,               --      sink.ready
			sink_channel       => id_router_001_src_channel,             --          .channel
			sink_data          => id_router_001_src_data,                --          .data
			sink_startofpacket => id_router_001_src_startofpacket,       --          .startofpacket
			sink_endofpacket   => id_router_001_src_endofpacket,         --          .endofpacket
			sink_valid(0)      => id_router_001_src_valid,               --          .valid
			src0_ready         => rsp_xbar_demux_001_src0_ready,         --      src0.ready
			src0_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			src0_data          => rsp_xbar_demux_001_src0_data,          --          .data
			src0_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			src0_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			src0_endofpacket   => rsp_xbar_demux_001_src0_endofpacket,   --          .endofpacket
			src1_ready         => rsp_xbar_demux_001_src1_ready,         --      src1.ready
			src1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			src1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			src1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			src1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			src1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux : component HostSystem_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_src_ready,                --       src.ready
			src_valid           => rsp_xbar_mux_src_valid,                --          .valid
			src_data            => rsp_xbar_mux_src_data,                 --          .data
			src_channel         => rsp_xbar_mux_src_channel,              --          .channel
			src_startofpacket   => rsp_xbar_mux_src_startofpacket,        --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_src_endofpacket,          --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src0_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src0_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src0_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src0_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src0_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src0_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src0_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src0_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src0_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src0_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src0_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src0_endofpacket    --          .endofpacket
		);

	rsp_xbar_mux_001 : component HostSystem_rsp_xbar_mux
		port map (
			clk                 => clk_clk,                               --       clk.clk
			reset               => rst_controller_reset_out_reset,        -- clk_reset.reset
			src_ready           => rsp_xbar_mux_001_src_ready,            --       src.ready
			src_valid           => rsp_xbar_mux_001_src_valid,            --          .valid
			src_data            => rsp_xbar_mux_001_src_data,             --          .data
			src_channel         => rsp_xbar_mux_001_src_channel,          --          .channel
			src_startofpacket   => rsp_xbar_mux_001_src_startofpacket,    --          .startofpacket
			src_endofpacket     => rsp_xbar_mux_001_src_endofpacket,      --          .endofpacket
			sink0_ready         => rsp_xbar_demux_src1_ready,             --     sink0.ready
			sink0_valid         => rsp_xbar_demux_src1_valid,             --          .valid
			sink0_channel       => rsp_xbar_demux_src1_channel,           --          .channel
			sink0_data          => rsp_xbar_demux_src1_data,              --          .data
			sink0_startofpacket => rsp_xbar_demux_src1_startofpacket,     --          .startofpacket
			sink0_endofpacket   => rsp_xbar_demux_src1_endofpacket,       --          .endofpacket
			sink1_ready         => rsp_xbar_demux_001_src1_ready,         --     sink1.ready
			sink1_valid         => rsp_xbar_demux_001_src1_valid,         --          .valid
			sink1_channel       => rsp_xbar_demux_001_src1_channel,       --          .channel
			sink1_data          => rsp_xbar_demux_001_src1_data,          --          .data
			sink1_startofpacket => rsp_xbar_demux_001_src1_startofpacket, --          .startofpacket
			sink1_endofpacket   => rsp_xbar_demux_001_src1_endofpacket    --          .endofpacket
		);

	width_adapter : component hostsystem_width_adapter
		generic map (
			IN_PKT_ADDR_H                 => 49,
			IN_PKT_ADDR_L                 => 36,
			IN_PKT_DATA_H                 => 31,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 35,
			IN_PKT_BYTEEN_L               => 32,
			IN_PKT_BYTE_CNT_H             => 59,
			IN_PKT_BYTE_CNT_L             => 56,
			IN_PKT_TRANS_COMPRESSED_READ  => 50,
			IN_PKT_BURSTWRAP_H            => 62,
			IN_PKT_BURSTWRAP_L            => 60,
			IN_PKT_BURST_SIZE_H           => 65,
			IN_PKT_BURST_SIZE_L           => 63,
			IN_PKT_RESPONSE_STATUS_H      => 83,
			IN_PKT_RESPONSE_STATUS_L      => 82,
			IN_PKT_TRANS_EXCLUSIVE        => 55,
			IN_PKT_BURST_TYPE_H           => 67,
			IN_PKT_BURST_TYPE_L           => 66,
			IN_ST_DATA_W                  => 84,
			OUT_PKT_ADDR_H                => 85,
			OUT_PKT_ADDR_L                => 72,
			OUT_PKT_DATA_H                => 63,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 71,
			OUT_PKT_BYTEEN_L              => 64,
			OUT_PKT_BYTE_CNT_H            => 95,
			OUT_PKT_BYTE_CNT_L            => 92,
			OUT_PKT_TRANS_COMPRESSED_READ => 86,
			OUT_PKT_BURST_SIZE_H          => 101,
			OUT_PKT_BURST_SIZE_L          => 99,
			OUT_PKT_RESPONSE_STATUS_H     => 119,
			OUT_PKT_RESPONSE_STATUS_L     => 118,
			OUT_PKT_TRANS_EXCLUSIVE       => 91,
			OUT_PKT_BURST_TYPE_H          => 103,
			OUT_PKT_BURST_TYPE_L          => 102,
			OUT_ST_DATA_W                 => 120,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 0,
			RESPONSE_PATH                 => 0
		)
		port map (
			clk                  => clk_clk,                         --       clk.clk
			reset                => rst_controller_reset_out_reset,  -- clk_reset.reset
			in_valid             => cmd_xbar_mux_src_valid,          --      sink.valid
			in_channel           => cmd_xbar_mux_src_channel,        --          .channel
			in_startofpacket     => cmd_xbar_mux_src_startofpacket,  --          .startofpacket
			in_endofpacket       => cmd_xbar_mux_src_endofpacket,    --          .endofpacket
			in_ready             => cmd_xbar_mux_src_ready,          --          .ready
			in_data              => cmd_xbar_mux_src_data,           --          .data
			out_endofpacket      => width_adapter_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_src_data,          --          .data
			out_channel          => width_adapter_src_channel,       --          .channel
			out_valid            => width_adapter_src_valid,         --          .valid
			out_ready            => width_adapter_src_ready,         --          .ready
			out_startofpacket    => width_adapter_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                            -- (terminated)
		);

	width_adapter_001 : component hostsystem_width_adapter_001
		generic map (
			IN_PKT_ADDR_H                 => 85,
			IN_PKT_ADDR_L                 => 72,
			IN_PKT_DATA_H                 => 63,
			IN_PKT_DATA_L                 => 0,
			IN_PKT_BYTEEN_H               => 71,
			IN_PKT_BYTEEN_L               => 64,
			IN_PKT_BYTE_CNT_H             => 95,
			IN_PKT_BYTE_CNT_L             => 92,
			IN_PKT_TRANS_COMPRESSED_READ  => 86,
			IN_PKT_BURSTWRAP_H            => 98,
			IN_PKT_BURSTWRAP_L            => 96,
			IN_PKT_BURST_SIZE_H           => 101,
			IN_PKT_BURST_SIZE_L           => 99,
			IN_PKT_RESPONSE_STATUS_H      => 119,
			IN_PKT_RESPONSE_STATUS_L      => 118,
			IN_PKT_TRANS_EXCLUSIVE        => 91,
			IN_PKT_BURST_TYPE_H           => 103,
			IN_PKT_BURST_TYPE_L           => 102,
			IN_ST_DATA_W                  => 120,
			OUT_PKT_ADDR_H                => 49,
			OUT_PKT_ADDR_L                => 36,
			OUT_PKT_DATA_H                => 31,
			OUT_PKT_DATA_L                => 0,
			OUT_PKT_BYTEEN_H              => 35,
			OUT_PKT_BYTEEN_L              => 32,
			OUT_PKT_BYTE_CNT_H            => 59,
			OUT_PKT_BYTE_CNT_L            => 56,
			OUT_PKT_TRANS_COMPRESSED_READ => 50,
			OUT_PKT_BURST_SIZE_H          => 65,
			OUT_PKT_BURST_SIZE_L          => 63,
			OUT_PKT_RESPONSE_STATUS_H     => 83,
			OUT_PKT_RESPONSE_STATUS_L     => 82,
			OUT_PKT_TRANS_EXCLUSIVE       => 55,
			OUT_PKT_BURST_TYPE_H          => 67,
			OUT_PKT_BURST_TYPE_L          => 66,
			OUT_ST_DATA_W                 => 84,
			ST_CHANNEL_W                  => 2,
			OPTIMIZE_FOR_RSP              => 1,
			RESPONSE_PATH                 => 1
		)
		port map (
			clk                  => clk_clk,                             --       clk.clk
			reset                => rst_controller_reset_out_reset,      -- clk_reset.reset
			in_valid             => id_router_src_valid,                 --      sink.valid
			in_channel           => id_router_src_channel,               --          .channel
			in_startofpacket     => id_router_src_startofpacket,         --          .startofpacket
			in_endofpacket       => id_router_src_endofpacket,           --          .endofpacket
			in_ready             => id_router_src_ready,                 --          .ready
			in_data              => id_router_src_data,                  --          .data
			out_endofpacket      => width_adapter_001_src_endofpacket,   --       src.endofpacket
			out_data             => width_adapter_001_src_data,          --          .data
			out_channel          => width_adapter_001_src_channel,       --          .channel
			out_valid            => width_adapter_001_src_valid,         --          .valid
			out_ready            => width_adapter_001_src_ready,         --          .ready
			out_startofpacket    => width_adapter_001_src_startofpacket, --          .startofpacket
			in_command_size_data => "000"                                -- (terminated)
		);

	irq_mapper : component HostSystem_irq_mapper
		port map (
			clk        => clk_clk,                        --       clk.clk
			reset      => rst_controller_reset_out_reset, -- clk_reset.reset
			sender_irq => cpu_d_irq_irq                   --    sender.irq
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of HostSystem
