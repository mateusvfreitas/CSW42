`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ng7z5mwI6mQRllUEyprRk0wiTnzc845VwG3yV+s6pIxZB0oy5WiOqZQIWuNXqKdK
k/G3tMIuw7zjlgtpXXktBtvTExxEgFDlXs69MniBPChAYEZNW+lJ9ug2ZQsI4d62
haUwMIqZvQvPGv5O4dovVG5yXhLDFYoZbEfmB9Y7pmwcLAita/mPiI3vtFjnAEz/
AD2hRgqVwKESl7ncSeGUApha9DZll5CxCT3x/yycwn24XeWfqH8aAecKmZpu48p0
zSo/7pSbFA35gR8nuuSvLQ19VmzDYPRrzLVrsFkmPAja+pyBtL+na0CAgVBr+HH0
P80a60c/nGXY1DuzUlBBhTEYJXssK5eVrWenMplzWcdc7aQunFxVhe7xdMOL5NvU
dG0y8MnpNAQUaQjnkroZ0zS7+rsYKfvcoEC6S7gbwyeHHbemN1bNMc0SoH2ZDO6V
PkHUeqi1NKeKXdh+kG6s9YkDRdVYh4tgfkwL7a6HTYHvkF9H6STBSaWLXZMaAskU
QwX7IPRvZnbNb+XLpEEmmWCc8l5CUL32Gz5PAMZdgaXlZlto67CIN3P0Va3HXZFy
6hPuIqhzVF2cns+PRHUe4GlY379vt5WpDOLhelXVXKdgfH6h3D+OYKdpaVmRbOH1
1czJ5xwaWJqtFkGkX8ET82OUHj/SG79NStPhet7RcsmG5nYIPz9ThAh+Ii+/98LL
WEhYpuS1iiwfRGIEEc8rsj4+iPdNVlA//OVSDeMmhsP3bNLB7CbQD9mPj0uphuWM
NyWKBXDH1S2OgIrtqneH9g8cC4KhYoJYpqZFSw3b+eWtK8I0eVbZ5FKN8psnvvop
TdSnsn/kCjNzs/WaF49Met48pv4se+2D03ICNUGREVF1d2qfYYypcXGe2Wj341oI
MqononWTwB/YSdMgZxZK1BY6zWQFQtD1HsmS5eRXtwwpFOPsIZgWw/XpmlXDc4e+
I/kv79TGjwn1S5wuYWuMlXOggtGz9NqUN5H/i8aENQ/55LzW4Z7XdFClRQvyvqhw
L6o3a5dTA/WJtF+6+VEt6u+0wiqhb2weFg+tX6Mey/pPNvDuxRe3sMtg7bOu/PB1
XNFbCSJuiZNv5xSpKE40RkMOQNDSnbQFhwoJPw4dApMo8eTTgIsC3S+KiK/pFuDP
crq+PgZfRdbCfYtyL0yo1w3eV1MfNAZQmT8UGFqXKYirINPQJ0MyowM/4U5/p121
835TpKtFbVwXC6A0o4q0V4hzaVYG9QV8+3vtqIQCFfQ4MECC9vZDMz3X0Pz5nOm1
BbPubqde74FzwrKqpbRiBSeqsL5UJxsB64CYpE5Z/yTAM+O4c7iKBRuLbxqdqj1l
/JkMhJ8MD8uasTcTyoCdzqOKUcKNk4sEdgKiRaIw9DmvOHasTOt7o3F2l8R2VYLw
+ydqTEw6IGGYM4a2aFA61j98Y5ciF9JZEsg5ON4tx90jjsKJLNsrcCPw8qs18PQH
DhPoS8F81ASHEePON5rb/oEqOyKqhPGOJdlfrTlXb+gr0Gw6yOYSTSH4JUQ6Dzg2
UoJnlQl+M6mKUuj2V3b5TeSHGXHtH1VtHurIEchKaRRdEYpi2lrGk97t4cKujLFs
gB7oXYeR05uxACBqqyIPJziXq2fR1GgyadhjADU5/3/yG2/BG+q+zwQZuv51tPso
r7JvKd0NlqPPPQgUDReChrQ4ZpHeNAL4CSirpDMK5QLUmBMc7dRr5LhLgYIP9A3G
u1ABY1bbF4iErwmPGmRWdJsHW0Bq/Yc+4IBEC8pIijwoE48okZldZJTxcxfmTC8A
2VTnlzGsgUG0I3mIU+6QCWbHBnPifiwg/CYzPICQdY5z3qVKYLHOzHOmT49EMuPH
WZoG+rRP2OJ+ZwxhpCftcjUkgh2WbVmGd020eJYVOlWBUf0Lgy3LnIVk7/YGOQYD
p+W9+sYfN9uKcwz6IsnCFO2ljrvM/30Ed2N4k/C62Q0j3F4/ahJTaVSz+aYHUE0y
Bo+3Kdd702XNVOxKsFPaAi5PxuKapozbxz8OE8mqB46UGRq/G6lD0wzEi7hFqWN7
Ru586AcXb7fDVpsF52jtCfR85IRzl5nRld9WiF6rtZsPDO4wsq6S1jjPw7mE/N2G
Lfs6Jep5nnUkgAV3vPRhcarkpK8t9/LXQY4NEpcshmhwEY+7iSbg5yU1pgyNreIC
Xsn9/J4cTtI2Co8ObLx6MfnRZvnmYjhgjX0Mw0H9GhFSpjImbxorYl+qGfiJlmGj
jYAgqjAH0Lp9aTypyvbwQX7yHVrUtkf6PqTA/igyq1t3/fG+LjIx1BVvd9kW0uRg
DHAPNwKSBT+0BI18fGzMU9NMr6KqUqDfts2EByLTWXneS8SWKpvf1tO8JzuS9ipg
0kAa6J/xmNBVIkHvxAuQ878OMYQVBFHThqGlkJlxqaUrvI7jkBAyBVqqpTJm8AoX
4vB+sUoM+gO0qxiEBAPOR5dy33rwOn5is44NPKOYD9v8OKd0ymFnknrOgcSVoU1A
/Y3Bb6W8aGUXvldjD9d3iGrPHyGZutCPsFXaiNvzL87N8DsinItvGZROMiLHd/cO
Tz/kXNdmp9Q9lrSDgXQK3NfQL1neQWy8vHxvydNniTKClA9M48VfDFZ+1R45eBrv
PBK46r9QUrkZmCI4XqCnnZC2MnOxUkXRkxstr8Muq7NciRso/EeWm9wqIqWDOu/9
ma9sLwPKc64/kzPOP3HQvjApoga894/FQ4P8hmsz7F2yPD1bCle4gv8r1Iqdr9yp
9U5X3uvrJSFFwnnw3D7nz4kbts2tMN3DOFU+Fc6xsByhoez3mT0qjZ/t97Dc9jsa
1JCDNysF5wY8PnBM27KqQPwCv5INYNaHaVMK6OiGK1XThVV5flGjH0c0SrxH+DMM
kKe+RvD32aPk+YEIXzfE97fsHxojl5TFTUN12sgi4J3kTm2afMNXlbxcFWPSwS2h
iL19zURUr0r8ygXp6ImlI02PG8Jk3T00fibrzOuLQvIt+71lENbLw7PQyn3/CWrm
AbJQEHeKL/2IOx/Vj9WVWvD6F4Sy+Zg67gWsNhZsunC0TAfRxE3O88oec+FbrN70
indLg1qtqVECGMjhfdCEa6OtiCCOC/z9t3ZNqSn/b5uSv5ADImL0cEsPJTX51eQd
E7nnzCwu9MOAhKxUEUAbO03QSdgrMEG0stdo6m04DuwcbPr2ZOMW4rQPcOLzrxcM
WL9+vGcTLWFMCkz0/KA7zYP/fdY/iRo1GXfdtPsmNq/bD4M1XgiNJSxClqkPoYEa
zNMygOI4WFrnqWncYYE2mTAS+GaANhfRkIP5HgLMn6tG0NQpnzwMBKduukFRaZx4
Pao1AzgdZLn7T2omSyTJw0Q6wj0sB+cqhS0NmXylsZ9Ru0ID/fAn7dUJWyKZYDiu
xQVaV/uOEWPCHJAATxiurB0KUXJHGwgdu8+STDKLlZHSLtxChhNGlRatky9IV0Q8
50uBM+BHvGO4D76cBGuw5C3gl741cWHejJuLLfe3v8AF7VRqKEq2p1sXZJkO/pIO
VXG8cPbpKxHQiA/oNbzMHCPQKOGq+ceSX6rr3lexc36ZCPT7Jvhs4Mdqevh+QS08
V+k9UZ6hm1ZgbJL8nkRzys5sAOM9dTC4Nn9egQ8vW+yavGnEyIif+cT8l3YlGxUH
ki0aFCBdhFT5YYblatL7Eqsbu8tYX1hDdOK4Xnte7ouhJG4UQRV9gu9VcanVDpBO
JwlcjqBICdzuAQtdqtmw5XxpXj/9NXVvsunpBKcwsetMwKdS8XQ6/eau5mzzp0kL
8Tgv+oeRXSX33sAwzfwF9O0O7U9HeYOnszlBkgD2JGNaPMwbJpMZHjc5F+K0XzQM
MDdDOHnXfhvE8XED4yfwgwgH96mDWZ2pAGhs5zZN73TklDKth0fH8JoLb4ebCpxe
+hesviri5XYf6WFNa55MMrg+G9wtg61Cm8eYtn8t21MAomZJxVzjSkp7TR8DGZP3
EY8r+Q8bt4B170PeTEtWDcEd15zY/0oCfBr6dwmUy1Z5wpsJQGqcBOmu5KAd1nAa
xj5SWnyE7Z2phvAYcPB9Z38EdnquAEoVz+dHC+3sn8yEm9mnt7GcC7AIqpYoo7BL
TODV0o9s2JvMaaShQ8d3iChHDm1V52ujQfjrDZBGAD3ZDSqBIdj7q0HfDdBxgANC
ozudcDnUNU532jpxzPI5DW6IeTyufDTAYnEiFOi+SIvN/lLhXiLilf1fY8B09qTu
EGUDkGN1O7AHn25+UEjFGMbGmsW1TWG++5rxX5ARjl8DFqO8vhovms81A6PtmdMI
22M8COcwjZ+RQ7AVBxG6pHqmKQzyFuKlbvkQkUolimrWDRMkOTU5NVZzF+4by3nW
tFIk2/co+nVu8rRXzUjxK24CxbVn4u/FhhHUE2+Ydbxe+t7ZR5KrZ8+RjGZPysO7
MvN2K/7Af/ruuRdsR4Sy6JYhT9XBzW08bDMGp8YIt3P060v6p7BJtvsqki25lKvU
S3rycvwzenKrUsYvp+eeyqFwZRjXws1dhjYFVWVJWrzx9iA7/s1DoTWwjsW6IFLG
xnxtmpddAnT/ADPxU/1FOurY2AMHE6cT4iufVCrfLa+n1aK+9fCPV/u+mLAEtsNB
KO/Mar0/9dxJDbhO6Lvq1UzGcBNDIjBDV9/xoIuPFRePjG6FVrgrcMu7JKDQJZoe
dEwIiTrAlYhO8/7ZOraoQsU44RMgt0zpCbXT9IK5QWzX1rHIcIC/4/Iw991ya609
BUTL0M39FJ3waQMrGUWvZlqhBiHVPpDtSsSbJCPew/Q9AGg2GLm7itpejeepXXKC
rk188ZyY9zbwy+VrH9Q4Lnl8Xfi+3u3qVYiiAc9TpBfP/vfixaA30ET2XFqp3U56
fNv6KIbCwjeL7/eJKUKXHY/reBIQ53wqZ6xlaExq8eKDHbQexIdJKgVGV1XguihL
Q3z4Amb6FeYX1E1R/EHGUNoerBoiRAhDA32L1+fVY/rODM+mJbbnaTuoC0SY4K+6
HsswJ/3xcJS+kn00fxR/wKqvYf+0jJIt6OUk67BMuDOoXEVP+X0shPF6fRD+5t9k
Cj3MuDSXPkvkf0c2k4u7sVv5G1JG1Nq1bu4xPPB4LnsSPKOEab/tGyRdHc9hEk/J
BFbxe3/JnQk0y0hE0x6m2h7ibswMeeG1LcnyU8eM8imxitGeMemcwXyiKC9BcpXT
Xa1sRvffRarIFmr/BdMsQNl5rFsd8GaCJ8YTCU/S8Cv7Vv939EtgOvnBfpxoeRF9
aFRgYqwaDoaUuirGpaLeYABexxo8l5KAwjnpNLf1Zn0qnhomEjBJhKN0be4F6b4i
7P6LagNSmDH19BGehcwWN9Nze9R05vLkTpjqXcOBuVdwZ19OenH4dsMHeMlmTlaG
PS5A3tqrNgIgx7U/XRiLgvzdsqvvQDH0pAIAz4w6Xw6hepUbXl9O79LnVH5a59VZ
87SBkzXtoQTewgGufCwq+BaZNUt9AhLWNsbg0WXc8+kKphs+uH3yQXnQkJ7WpLNh
i/StpcvBNCIzl3KFjMkq2e9cxdjYPpysLe7IQI2txgPjkmvTgwIrre7SO1xCwPvT
dPF2me0xmS50tKjsgz613cH9kvrWOsqsN43ndiqfkeacpQVmUbLWpBxt8yxS77Xs
vWHqXhwL3VTThojvN3y+Cl2PT1QdhGtPYfZ4lqO6obGJDQ/4RsSb5O+n5SpmDbp4
5Lw9+mRBe2Z2ja31avTxHRxSS9OP7jd3wUrOPw/BbMCEUqojAScG+3Gg454TmbKr
kap7WhrP7JI/9g6MtXp3VaxzhSleP3F6FFdNFN+kSwnvnDn8MgGXFX2CzWlm6/jH
kyUVHIoII3KmkmTi3pAt4IUTb6jbHoqH03L4UZ0UuIKjqA/pbP5fZzTW4Cmjk8lY
V8tTBQGKdR2uuLUe8SCPH/QNVL3N34emQnelWbTjA2+RBKkH/FRRhaoWZFZDlJZC
Ncj2CcwNSYrAoIDsKhXxZQGbzpq8jFaFaR/sJ2e3rp9JcEYsWRNIBcxI7GIfKpRK
81EjAhQNUZ3kDZmQwnZ99R4kpH10sfLGLxbkMRDpZfSJhHszDGu8ffS+lrMr/o0M
QnYsB8+98B6pULHVHKctVh/A/3dEdiRNstNnoKbDBS3L4YgDofh6nI2PY2DuZI/R
RPQuKhkFVYCDfcReJ/UIl1p2zxSXMBRxf+lKq0zOmmQjbDe5ZKkzotJNFAIBXHO7
0KDp5/s7Aesgh+YwX4ExnONHJ57cPkLHc2sbcGgj1TKm184np4dt9t85WoYExMMR
FKNUILVdKOIn467sGy5/sjEee1DVlVCeWI10qimGhCHbP46Oh0OZS8LsZSiLwpYJ
e1AWXgqSpmEOdGkBBWeT7ZUOe8Of9byTVC87PZ+4IHWwuTUMUCO8JJaqAKDF6tfU
J5BaGQTJDVR+JwhFUY/OYprsoRFXJuNjRZU5D7Tk9MLoo4myWOpzQI3XVwHdT5+u
Ng4ktK/rL+n7gf1VRROuL6m8rPqwr1yZ5c37P2jPOO3z0wZV6MuCuO7kFUws9yAk
+f5m9F/SexQgOr+xnPK51iaLqWpm3nCIKqo+ejhflD6xs5+J4XzWGB+RGTMhd1Gz
FFHFhmEDaMGufzwEJyxY7a1tFO7h0laU3VJaWsvPdfews2shooU2Kz37P0Mzc7wp
vJZ4LfKhPKZ4DcfuSim3XfbkUZtWcvto/7ITYO5fnBBZslcxnu01tND9tCJBEZJ0
9cJa7GpVFARG3sOkpS7DHGtI3d61aBOtBbYR4qUYDNP4pvOjzmjILZEJ+qd4nu44
iU0cxaVaGXnYmwovpt/Lr7wleq/EauRhMnACyFZHrzeNHtFVCVwtfVBBarDdRW+F
d2smTLtmhv+d5sexqJWxM0UI8yVcDFHjMaiPU7O5Gr7qHPNWb3LblsKmoVKFt1Ef
/X/RJi76TDixVbAywZfR0wLECsZQknvw7h/+NuLypEXVEOMheG/3jgmvi47SFJcK
824qPWFXrknC0TBTS9WqP4HSwb1BsUG9aI5eeE+9UVfM1MqjXulaiVE4+KZwMTKg
riQ7Cbfzs/T/v8yRoBXq6z/KSEXMJSp5pCatrzME0xdAnikH9jgNht5+QRCUogmH
+gKcJdDP8LwtIiDT2/wi4WNcRYajf8ySu9M4Ilg2vvbcxVE2iXiyui2blMyAUG6e
7UbgSn3VyvA5XoNqGWjUnHvX565GfNuKLCNQx9628FJQi58Xje7qhr5AXkmPUiFK
YAsfn5mRf6lVHz0LFuzURQvRmrcw/mkTHxkuWekMJjN75O45j5gxMWI0gLCBnOmb
fRs+l11mkgkY21WlbCaldFNp3UwSix1sBd1R8sdNwSZf3r6n1a/9XmA3ROBHsjZG
0DIrIGzhwsUm/nddrtlXQDX0lHO99fKLH6WVLRJX8PtD6bIznAcxHLv4SKJse/PI
7PirtIZB3WP6m8YUCVNR/HqCpUrLn0eJSel+D2imz1NOtiXDLEgWCUW2C7lHP+7v
pt+9IUSop7gTaZNqeV18Kna3GCcNA9ZpAm4T6maPOgedU73QG0nAjwnX58fmKZEd
xMI9R3EgmaVIHvt/g7a4KTp+HasFtO17phywXfPKeQGMZqfc1es9mw4WxN2+tpYx
i7CFXHPdqvi5xwNUMeZZNEzN6GsZXztwTU1rAVvbFku6F8DUmufpRDux68eLD4cs
`protect END_PROTECTED
