`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
C4FTU74rk28ijaFMDEGMkkbOZeOnlorweG9h6fkJMojl0/P2n2NMKikGFN34Jeo8
lO+3M0QpjA7kj0ZcNL3oOcRVysc1PWEvZzAPzDdai71EPFc4L0vVy/lptZLUjpM2
Gkv28a7YO7khkJa4jOIjIkflAmhZx3Q36izDwzl5yzib7RxD4ufTRvcTGjZWsptz
sfdyOf0qBMMom2fJUxKKx8k+lbi30kGU1xNXd9KqoJmM+WConkVfQNVDsVEQKIID
fD1NDyLf/Xz4Kn7FgXLnhRhM2DNpujxmnERl3C2g6urcYtQ9p5yN3em2kE98fQqZ
0GCzUdaciZ1D6TchX1vZ2olOY0dD0iGn+IO/NQLP9V9jxaFmkwJMWUpypsjeN/Q3
7Rpk0ap+d49vDt0E7NuyGSmtnetQOQ3KPD0k9twa0ADp/UAI2IqK2xabHtT+oNnn
QFtd6kWO/0mmY1OHWl2tW5sm8UEBLEfxuFOcGVsc5iK4SKb2aYsIh67po0TIUg25
kF/Jog4+AppsJk0HZv9id7TQlgz59FbA15zjjYoE9HSpBZ7F8d+ofDcGv+KIRC8O
/Qz7CDhZLPfJYSz61Ls8UhKwn4KVkhYZoytJRuoxqmBncZiLJYyr6cXZr1FTDUus
ZkahBhCxmgODeYKlVUM/AcT2v392q6KJjGMVNqVAUxtw1x9RSg9NgaBDXWU1KoVd
al8F+Mz9tT1qzoGNyiPdnV42OVWyZfwn8Lgd2ZLuHon5A8lv8/1QfIMfY3gMidG9
39KNU8rN8TgyP0SGC/NKxpzYhqz6TvJYVE/j7ItDEnVIW+BvrxRPsZUX7RJM/sfs
WMBsh+9JWUqbcJu2HDfAhnbOXTYAQsJhqoeowtsbUZ3yRnMQWYyMCaj+R22xvxac
1x1UDQ+ARVeUlKhVJTdy7pWfUkHRv2hm75r4HFvjn+3R6a4SLZ3y43XxVyriCZKo
IRPSrbL57yw3ED3PQYQaJTYPXa9ds7kqWrK95x/vmL3FAvemsiqOnc1Iyhmg51EQ
kPBBHsECEYfm61/duSn09HaL+ZjbpU5M2UbKk3pkmREBsX2PTYaQ2eHiB/lGjsai
J58eAxr40FJYuU7O6Di6DZq4JJSlLLD0jJ04RfF/9oF2l+7A6kJ2p7OmAnDhEnKD
Q7UPUNfBS9tJSWvXoo3cSmTtUzkeTdmMwrusXAGeMgndK0HxfFHmNI8PW9ByPIeJ
rB5m91GmAzL6/JoihLP8e8hKmYC6FDzBCuEXAy0v7cOaBYbatTFJhqE8vSgEL4Wi
iI9dKDh/GQK7bK+sZ87U8LqOMAC5HDDTOI5UjnfpiKh9FgYu+DMQF9ogBK3y0Kq0
KgWbTUd/9tTks+VZZkbYSJK9FlMGeIzqoRrGYh6azRIJdXSsJObpHlBNmdtqyIbk
U4aEGwbnPuWbtG5hLgTTA9kTl824DncJitog/kE48iPTTqepNnKQemKD8cJDuXuH
8UB6WlCz5lyVcKkP42fns0gdg7+HC2L7KDVQ3x4E03hwCPMnhabRiqqAZVzD7qQ7
AqTlVwdBeX/nl1X12eawO5DYamcdqZyl7WcSkbWrjEZEaPuFsYyTukhIB9wPPGaj
L/dMz8cgYlS3V1H/+ZCkBsjEMuLKEAfl250Gn1Sax3L3BvU6RZk18TTinP0i0w85
iRQJh0sK2VW6eQe+pQBL7WJLQDx26ZF3IOOlmdSeQBL0tc4NQhdXF72StgdWN9ay
jF7PXMpGX0b/wwtDxwJpIRZ10nPNpEom8W3LiXsojof+J1AzUfKzAJVPF/Mmpijz
iOmhgZje+g0zk7e+X244gOHyLSmA4ZYpWB3y9zFy9rFNazt+thUrZxESvl/MVhdt
D2wU9IrS30fvRRuX8VBHJDS+dOyGVkc/dStwPKxXTI3dW7MLFK5TcqX8+6gbV8HD
cRN/lUW+horY5R+qORavAXL7p5ARRwauAXgAaRjypX6acQgusyOdMoCbN2Tce0zI
I545kIHkOqFdH1dvN9jON146l/VMerXnlpojuw1c+2/rteKeGXAjTYakMe554Nwy
HUETAdHJylint7jErRQ2RuNB+o0zpZjhuMHNgl2cyTe0gARYjKY6zXtcvQMJ0HgY
4iLa25Ufeti//rT/FEY2Nv6efBBrsApzS1ZTLvg1vmB9Q+AIfA7RRekCe+MMi5YQ
myNsy2yVgMy7/tYITohBI4yFWCy7PGIWltrWLj9UV+rhU/OVj44eG4Iq+uUWDLfV
ZhvGABOvB2F8/2KTy4PgkQ==
`protect END_PROTECTED
