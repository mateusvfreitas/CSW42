`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
t2VJo3S92X6VuMHKbu1iOXsIrX2oj4T7pY96CAApMaNBO7+gc5KyY1qF5hQq/9g4
L/YYzJAOQ37kD3txkYZdtyv8YCvzzq/ZtM7k68loVlJACy+MAdNIgyUdyHP7bICP
eW8nYNMu+JVbQyMjLdOvD4n8dI4VHavd7OsVDTa3JfrSIQP6tRN8QUFD8HpPmpP4
2TPxagd29xebUTztAzJ7zj6RNNu//bHer9ir6aHl9YnVV9Q3xljFYmddE+r1qe6b
tIJeyFx6tF/WvNQAwWG6iNEaWDtEwLvhfrRyD1AzjG86EKfbisk4uS5/hmzjydag
9W2UMM/Ml+KwImueTrjT21PMMLOnAS59bSd5HsmAt9dZDhvMTlgNHHprtgaqKXdV
JR0deRuxrAuSSso8MWqzE5ZwUDwyPpZR3gmwnzoKDHuuUv1/+yiG2qz8u8hXXOHH
/z+PxBs0BqsXM+x+uZi0M7gr9IfRaJxoVDFeC7oJz570TDzYeiR0jbC2rp8c9Lc2
z679WYsdufD8zvyaonNnxM420nU4fqyy7793BVsYHopCVSUTzy4tX/o28mVNAdyA
9XTJbjpLEok0piFSbeJwYiqyDYoP+NeTbcHeWuil0/WsowrMf3HbLYPg3QATWgVf
AQ5dZ8nXSZYl9VIy9eA3XrdZWFKnWbAarkJNVBdrhmdCY8J87+d0ec9oATiDlXDH
AkJZ/aiiEIglndkg3o+CUO0YxeOjjMbhJtx3g3XSCrqnvb+NmpOWpN5FNCI5dz0m
rm73H+accHV4qbjLwl7HObuXS5+abnqTH6QNbZBV4NwS6aMjMVLLg9CVOKb05Lgl
ErDoddPdiKLui6A2yWshDuvpCujdcW1XoXlYpepubyXQDMNlIKEBcCxCSCWwCW+q
lgXcaq/YJ8N2H+C4tg/iURynhMzuH2U6nAu8s7FhBYnUzUtoOQ6CZYQTcl5nzBwR
KQ/7Aimshg/xu7wSiBCxAUy+R5C9gaReb0WqoQ7z8xPtpOa9OyjNSzAtQuz4Bd3C
BDJxafHc5KHIbjUDDSm48sofPGP4JV+YUPabL38SRCMVhNzw5vzPQsZ6+eaLdLif
4ohRjFCqqygU49vOxAHtKroLACli++TBEXt5GdSQj302ZeCEkLbBav5TikJbw3ks
ChW8JDcaLlAH1n+7sAlVzP6gm13Jkt2JgFb1g2tFLHX5mZLptKONdZnbqiqmW2HU
cfGUHZz/TClrqbQbcj2VBQu/QNNl9I7/B40iMN32FpvtHD9GGJ6iz8muS1c6Cg0n
+Wuywg/UU7SdgkHyAXQ/r6p6R4evwOHnlD29ufVSc/JyVeIOUhH9K/4inbY/jOxh
Vuqfwoubfcev21wrZXqZxDB4wzaQOij0RW3cN/GOiHfzW2/lwDTAQuJwGro/wyPf
jrq3/bKp4ShguBR6Mdx6ktcXPZ5uYkTa1JznIfKDal2oB2YxpRwV9gpPpX60eSng
nzcbda+R9ZYFOsARwTTdaiVq4+pNQjvAo+T0CD11eVsV02yatyFETTK7xqPznfl9
5UR0QwMsrVrzFdftSKwmLKMeTR6cgowMESuoNcimDzxtlLRVQS4ikAkM4akalKWn
/sdPCQdVpM0wUxfLyYkl00wH9TFe3X2mfdYMrKFy3gDwmY5Gk82xV5Wz3CXoCIpR
y0dQOYhqz+xnVtHcsO4wkHDkv1b2rkRU8jn7hazNQbGoWDzjCbz8Pzm+MsxzEjxW
/z97+qCUZChBh2I4ttCfcwgXf73BVvR+0Muoo0uvmx1RX+UY3M6rQarPoCkGzYr3
Fh7Wnk0C0O++SwKMJsNmQQPQMux0aYkkdxnGS5B67kdu002D772DMeH3qWi8LENa
zbeoVgGQED1hXhqKhpIjUPjoL60zYB+Xcxj0hcsSz1wvHMXi6VP8YtRicfo9nggW
u7qbJzQUyV6C1coidp2xDtHWgchq8d/1NKo1cPvRYJ3Gjz43tTZxYLQkLe63j+kL
QDIlAFlGX37h50Tl6VQQ3jTgEBw+1Ta1tEPyif6xyaQ6ywsitk3CozZYhJX0SoqV
Q6I7eXHzsxkMS2iAZnb7zwaWY57oafF08i6nXXlZ7ZTtyUJLTxBQvpswcAjnAQEx
kx6QXVrVvvgKEN/wVQQacYJfaGFPoaBz9apTHC8QCBImBseQ8Cq456GS5cn78r/3
nfuToRSkmfCOK+4LlxdjI3lXSLMhZRFoJCKRKuW6/+9K8eTFiLsM5mr0+WGysLaD
GpuKJyGk1rfzV3Q+D0CkaQ==
`protect END_PROTECTED
