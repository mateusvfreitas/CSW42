`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
smpPhzMAUZGqyEbO3rJ2YVXfmoephXh5nC0bPoIQXN14TixS56BO1zQzcovTi+fG
5AnaWV6QQ2v+kbNZxpnlKAR2wM8W7WPXiM6EX3UQt+nwQJ/HhL9gvxh+1pLfpZOK
7s/g7p1aGtnDFOLudIfRDdvFfMKlAczDtJkscFPhFXHDwn4gXbrptVWE4/aAHb+a
XdH3EtjNA0tJdQk4afR61ub1NLAX0b0dccu0NpIjCvqBKO2iwzwt+HJNDIflXhby
By1xyQ2LepD6tyKf7M4yXytQjpFwCqIyOl3rfw3E7riQbBiiYpqD+AH0id9NT4X0
LYe9UkbWboRIqnjZGs+1QK0FW3xI1DriZGr4guXyI4G/BLHLCDobsjGne1ibaze/
kofieQNJg9/eI7mrySf51O9ljFBZjgfi8QtbKX56cJzvovWvoNlxiWP3v3ttbo8J
9mObBhiJ94nHdxsoWjzFuM9iLn9gyW17iFs495sK7tzhjMAWx4ggy9jRb7Ba5pGb
gz9uPDNeObzyzanR9/49UYq7wDuDkfyoaL7I44lw75Jy16eq1+1Q3wEg7rN0rf+N
F7WyFVBJchUcPrhzxCFtKlY/GIgOj6AcbD79oEqkk9TaHlv4U1pJSR5ZjvI+RsSg
iRDMriudyDRtizxS4LyXEXqyIzfKD1BeUEhO5XsaTHhbTRKW+c3V3eKXZYhmjLJF
mEeFFpeeukiyOXyineizozJ+c22z+FCF5Et1ME/+cr2yFWlRZlJq6dHoR3HPB3lT
ahjV0TD2Lyn8Q09x4+SvrsZvTIkmRmF2YeBNGPkqxbtwG0wM/SEuXivC6otEuNEA
+yVQejfN+EPdDu/JJBUYSgWS8oO4wtNSd54kx+XtQ6yFWWYMuIF9CC+S0/2itupd
qRDscQgLHMaJNcYgJuxY3If0B+g62y7bBMV6JRm+0yJJbGvzhrIUF+9XuHW7GD5o
2P7rHZd+a81RHRB6aLCQCVvTayCR1P6Y2dNvSijS36wGJxz9apRdtiZFNxXSpqp8
Q+LRx6a5FstUfQC55SZx/N0B4DmdZKzwkadG6UQTuBtgfrSu2qffUZLdGqulZXBb
Y8U5PCBvIgCimGWF2MsVjF6CFiiHTNNv90SfkLD4Rodg6l5R+PlBWYDHa7UJIukw
VfEFiZlDoe3+/GMU4VbEUQqOAQ4AkCY0o3jT6Si1kvdW/3xACEVR78vAOc5UJ5yy
muse4tS5ZjY+GccOZdajyCz0Vpw7lnhMizZFO6U3RbrtxX1OzafqwL4EQcjjWQez
aj64ZmRikpI0CwWTy0SKzhZQT8vuq/jXCuzc8p2PpSWWp+ynQklPTygIg1jJTfeB
zXzb46AeVqChDb0Pe8I3GWKrtMxzG3K3ugcjKw3eTJXO8b7Jg/1o2idhYDeI+MiO
UbK+etcgmfUkkjm+NnfTOFIm+9xxGtsaMNunaGufLqDJekXq8zJReHNPBUOeFjKY
0YbKClAglOw/hpofF6ICqCbHyXIXIZWpH9a6id3E2brM//FH4ve4swpTbJMKrUJW
SJP8nZGxxg88+z3SCdCEkTR/gM/atiGn4Dn1M3YUVoQqMIM29gKH3V7pI1LNoXQU
2Og5XXh6LNeLJodXoNlOK4Lo8JFloDW4MR+nq3IUpaRB9eEY7HiNwW5jl8fppdlK
1E0roUU6xAriLjAnpViRS+wRBWVM8WTLrppUjw0l1KJGCpf3qKqJjy7thZqXFF5c
teWLpuIvGhEggL6Rc1GRtvHMdX2BF+OnTvlpePkByqKM6FDH1R1weUTPcQ9tvUXK
0sA8uTbs1B5xic7L81FHF0ivClC2SrH55fL1aS9vOYPzAmFepfByr+0TOBCfmPg+
m/i2a0NdfaR+higIWwURWD4AJS8/QQThc4yspg/eh9Rt+2UL8kxLZChg6go5/qbB
bVGtI/fLtgPn3J87UcH7CDAEtL9cZnFOP6WnieSOC3nEPVoahXSRKzX3PV0GzodQ
ywwD7IeRd0yapIaDgrnRTQhvNKsvo+MohULS8VCS1kxwruapYf4ftTV6PXDdwNBz
UXFa0uCdzLkT1GY/O3DbM0+BBJO5pgBliIoR4KKAGdFzmgjj+xyDm9OHT/P4kSRc
wbCKCJxB6Lwj3pfcecTot+9YkW2uL2jXGO9Dx93bNo/C20AlnWXYa7r7LnlNLn/K
fGnLNggCb6TlvbYiz/GA+EK0sssVHR7mNdwQPl63flFHy0c6Aud49TWYTcg9QJnj
gSqbnJwvhlytuewU2ppqHA==
`protect END_PROTECTED
