`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TYbmATtOdIoduvmPOH+fPBCpIdVNkh/jcZyRbEoUkZRfX9HEmHY8ZAWpdPrp/FoT
ZDCdsWLrRj2KuiVPRRHaIpbaaaIEtvDqtbPnxkTHUnMKEagcZP1qxc4jmCbCNyaT
lfDio+TvkvscWKPOw4b2+NbkZPZaegVrNk7qVBu3AM8/zZpetcewy0bZhMvwj7k9
QhGwctrLSFiWlTxUV619L+zqLkWgoDgXRhrwHriIkf/wJ4hYR0fOw59vZSdDiLCC
AKqHf3Hlgsw3URrpBEFhZi4wXv4vvZqbTqDxlgm5K3AgjpPz6M6MA2QsNuDrmDhh
ltvVq1/4WPjb09iIqNjyQH9sWZ0yOn0SzYJUSMtFEt/jF3oIbcQBEk8Wb0fkJGGd
OS6H8Bu+j2IjBSrB+2VmpIXI4ZJJHQqc8Msv7lVkQML9cnYQnnqOzezIqkTAGCYf
FdtklMz+mvkulEF8zRffgVJeP2DDrGdQKNpL1+NoIN0LxgDi/PnVgQU3ND1IWiti
A6/UwGl2aMqNbfvvG/qXVs0qodeSYCkr2d8EvdPcHIg+oFZmUOJokE8caH/fLiYN
GHBv8B3d18xZO7f0q5ASdyCxUdkDULM4wXVVwlD9ofnefDJqLLySrz/Ez+VyjsQq
YA0OTC/00orppx4KZCwBhIDrTTheSe/Idh9RCodtYZP6xRRc0H5BhYm/gKW6+LiC
BK6uMIHVCy4/U/wClLdeCp02IhwVBvDKdhqXqYuLfiMyfG3GSdGiqKS4fKMBEvPe
HNUG/uCVitDPXV9Kz+XrmvdXjRIWdSOqXg7D8OZSADZ/Nr6PF4Z8ahqyW+AG45xN
71QM9WbheWMerISOIIGZZDEdPXX2OLtWa1n4gajsG9xFT53ovhBSUryvmgfmxQ8t
Vzpl1fLqoZVBbyUk8CiZViUjkTRqaydIthZqTod3t5gygvh2bMF7I22iApdmlEJF
FLS923hI/UMvqLgy//KUxZPp+2w9cQ6UEvxdwxretCzUbbOIgUK+HuFt4n/pNQIV
go9QvQ0BNmvKt9jQ8tnz9msGUf1jMitNbtItlPPXB4wspOpMNUx8oj9vIBM83kBU
RA2LnBnvaJotTHmC5FM91CqNkkGfqWp0RPxxMRO8DVJAvb0iWg+VoPln0Yg0bABv
5oK8ViM09MmElHpQZCY/OgRutMm1hxDm1eBp/STG4Y1Q8aZE8558gEGtlvEs6j6q
KUHVU/iIrPt2QITjfyyzh0fgCsXTQ/lJkMsuJ/RRbGkg0GsOiC+f89IVkkU/SE/V
zlIp8X6bfhTSEYC/5/REP6NzSzN+8khfSi+qddbFEVQOdBUFIi8QfFfIUBnz0IV7
bj184Virt+VRaqeSU9HgU7Z7h8znUTeJHBjCU0phLlxkC+zS/0DsppXMltacb98y
ngfVPxcz/EYkqGfpdR+/W0pWLUrP04Rmu1Z8D4K5SUQroPTSQyFUy+NX3fvWkUa3
vwtZZuFt0Arbc+QHQne/djq/9b1bvzFVBJ7Z3w8XsZFZf6xXteWip47H0GNa10DF
fQ7ln/Z/wSPru8wB741bDQ0msSMfIw68Q+0xHYri8vl34LrdmpDw5DH0AcoqdPIb
gdU6BZeFrF4lugkjvP6Gh5HP+m9M2lMq+0B/3BS7kat+z4/HAwvTSBS7bRUyZvUk
/z4Tb7byMyfjgEAbr9GKgGaps/v8y9aBIT9lWRhNmWqQLhdohegOjLS4A2Z7S6w0
QJgGF1xkDSj0zMSWK3a4JACjvz0L4PKKX9wiF23QwjcGhrj3fer9ZdLjehpqsSD7
YunoH59/9AEvtXlak7iyU0QiyJpPmEseHb/CnvYCv0f7vOQtmT/BWmdaLtrqpiWX
6Owmd6H2E8rJj0ag0N9niHY6r+UPbafQ5vDrM0YQRwviNtPb9+TGi53RZRB66HsQ
d3lNqyYNbcTvxHy3DXthU45CkpAXdhRmpwFQEoljB3W9GvXTA+rSWfxKmr94rAJO
57gk8sbh2fSAuSUDZ+MuVA==
`protect END_PROTECTED
