`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dqgXNN6CQD9QVf9ZqWQsmNPCxCNUkOPCfX+llK397T72Di7cHeL6flR4BSAaEmNg
K5Qvr807Anho/K9KNAVNld7zZfOnbzzBb4lHrtUggvvuCaS+hn/x8MAugyD4ZurF
PtjK5CRexbfXeONlhz9pzI4X69XLAeCyhdmDEFMJkCvYGfvN5hFI9duSt91oppEF
VNUXlkJ5XlpEdxZhmXWcsFwHpzM6R66GBqLlNwKy6JBWkEr8ls48bWID+8EwRbIu
2Yd3ZLb2ZtRIq572HrLj6HvM/B4vNBwNmkOEF2l1gQRlFoQ72H1D5wqkigICIhuC
EiZWZ6HTLCV+ymPNP9XUZBtwYZ3mtWw/ujiIpAHiMDMm2O7uBujau+PnJFw9qHB/
kVSKmpzCyNRKeRbKkvV6vPtIVDepbSn0hME8Dw+rrVElyp7T1l1gWrzdagyPbd1a
tFuerYFv2EaAVYbHQuegeIGJCn0fNe1W4KaWCrQ51E+wO+iUc5OxZ9iRpL2hpX3x
o5SbuLM2yaJPYrMrYXtz2ohBknDANCw5pR9qpFFZgFiaEpA8WnFxkWpMoRY+Xrj+
HHqS+AJZRu0nJAkiPHNU/Nv9Uxolf98kPW3gf5pPmx4hXfw/2dngQ/EogsVVwHg+
K5fEOraEQkC226yFiRWgOKe9BV38lpdqV068/3jFsnlzd8/iuzVJAKHK1X8HVbJf
jG2wf1EoCZ/Uw3qt2aSZgDLOrgqdvvV2T6m5hD4C9EKlldsM+LvCEnZ3KE7oxJnS
XdcdMM2et4429YBsaXh1cgCCkZ15VyXpyaHlMTM1Ned35S6w80jhw16VxM7WeNgy
UnvSVe8/h2Ms2WuwjdpIGht4t3dpki1S5WPYvCRc9i9wTRUJ9PLW4KubQSRh9RRD
xTzCzz2C0OlowUhS2HYvsg3eu3YrMSTopkz5qrwWAkY2UZ7eQ+1GSX11+qia4urU
NoNfm8PyODOUIQ+UvI7wxVHRGMKcC/NN1Ck96p3f+oMgYlD67/F4VLmY1jshcbVo
6euxZGSgPT2g2GBwFNt40XuoXVa/wlDlYyWQB8rMGRphZCgvM0R+t243j236C/uR
zthXB5XI2dT/0T3XQaOuTwgdDFk069dafoqjznYt9LG/+WCtJyxngVLup4nw745q
ERMw7+ZQ0h3STOarNKP3QJst35JVIagE1lny+nEoNkstllVS0vYpx0MAI7C/KEjm
YBCfuB2jszdpWSD4BxFUcoJ2ptb9DseRZoD39ofCVGBLX8xvGS0jDr1WocEtkGWO
WPnXit5HhDt+c+x8EWAQi7Ba72fTTD02isSKkqomXnlgGODthsWbQAfj110DF5wm
4/rPqInLfV5MkrBhZGXbFKw/9pPEL45XuuP1O1ioBn+nOvmoF8q5DE49zrYbBb4m
tkWaW8ffNEg4u/q6dIq0kQUY706lWVf/ETcz+VR2ixHtYNuSiC+cPiqSeGWHrwUW
4SbI9fpd649xnngyWdOHeQAasvYUzUvIEAyggJz83vzXuVc6P3S0BrApGnZ1+27k
WsEqTlt7uVq+yGfSdHEyAY5JHrHZ5Kk9FmsTLZF0sbAh/gWRH/YMGWN8ri8zSJPD
zPJH9eEFIMjD3MPbOg1iNwvu/YG+MgGanpqrdUsn8s9Z41fAnNub1xswx0Lzb6eX
RDKOg1aWVeWeAm3XY1aWWO7yapp1o76/rtghYhOwSYljBUanYjnZNOBZ8sU1/v3C
7D2VEmu5qmTecQfS8+sYZPkvmeC8g9GwaPynmL1FFfb04400LalmrsrnmQtinnqs
KUcImmmLlbkayXlPsn3eMYJMsZv+yKFvGARXv4anYLx/t5ONiI2sD5NKXUB3KRLt
wRkXUHNxZUNSZerbMgizdZJsLF91/lTjWPkBbBD4+41w1yER5vUXxQLhA2WR9xYS
s6kQF5OPTGnHIdhiOIQ3rIzj6AxR0TREQzb5fQ24/BO0N2OOT9xtY9GpUBCKHYRZ
vrEPEw5K3HPxrQtDa/vOf1EUd8L0Jkf2WMr15w/vNkjrbYtd+R9bekTVWNveS0qi
`protect END_PROTECTED
