`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
jh5TopgQsA7fE9veIyVMQLRhzT1WZNuJw7SkiJdNr85ob2j/VslBxAhRDpykw0Ap
HrMMzzXSd1PmCtPdQVTEs1Q9cyS/JOQJqmL1cesfC/AeiPn/18nj3BwC4pAkn3tW
zIyk6aUbISHTTIlYGHp7Tb3OpjZsNvSaltOHqA7fUwqFwAdR+52/+wlaaxZbaebT
gvLEF4/T6S2DmzGJZ8qwHg3aEy/wU1E94+Sus6GO5cj7eIhGliwYpVspeYGs9qQs
O5U0bpV2lazEvpVXSiUCwgXLn4mi794yoV1TrOTNL+9QTOGvxpW5yRJraH6ZQrIm
/vePQZKC/o1UQ95zvyePpYRGIl5udy28OZ3KQGuv2naKVB3Xvk7bP9OQHDK6KFkm
V0vnB5wSSxCL5Kafjbo5orXXQCaGAbNXQRMyNqUdZJKmS7zvOtQIWoRMEON2X9Ez
zi9/Di7v27SZa62qNBGw+xQP2f2cHRItd7qQgu37kTHcx21SSUeZtv7b3tRiR843
URaYjkVdtg01zdhb/Rn2BTzZjj/9YJ4Um4YMwfkTzQbq71IzJQdEofD1b8T7H8LL
aIF0RSPjl6QgAFN5cWC5PMT2Ty4yEKfGV6NxplPZh5CzWlnIvbQAtOc5S0SLQUfB
R7aUJ3z0SNVyw1+96ZmeP+a1FIJ/Gj7f47DTRp20oOP23AL9bFoH4QKGrREkZvLa
Rixu3jX7afCt9bDpohz/pYlpikQWCE4Ep6h3JT9SICmFDAktFr9u3PUk8W9owx/k
bhxrYye4Zu7/bFUR8MJgByorVilGUx83WMw+IuXc8CQWSJ2IcTJSCCHccxKoabPV
YoxC+GsLk4IOvIYExE/+SfJVqcE1YGGUd8nC+C5EncoWgD8/h2d2JQ3OFy7EFzOL
eEJmZLtyh/k/5vlzH3HZqYaSfT4SWPZGIYSNB2Mh4QCQtfCWanSGj06f0hjD1TNd
qtbaiNfkqYSvde98e3PJ4dYe3PFi5YW5AvD282WeLD4nnvIWt/cm97ntyJuqCdRP
T0lIWRN+nEejDws3BHn/tL4MS++OMBCJSgglTYGxPO1G3Jo67dVGtLALtX2nLmg1
COVEFjK07aq+0nHBFRPBSH/RKLPPJLzymcP8iy8VzeJdcZYJrNZAKtnoStQ7pJSH
Y/pd21xHA3czJVspRAxBHpTii4RLMVTpkM9BlDgOM8CwKiFlEcpDS4LMV1FmPxhO
vB0C6Fy39eMb3k8ovFvw96RvZlVxFFv8kii0tMSihIuBVpt/1EALQXTjkqmije+l
XxegJSqpQliZKwcz0o9eRceBynAZKD+MRSbjVjKduAqeifAXZPv3HoGNnqSDHWRR
cYFO9T6i6jLnNo0h5itnY+zXCwvoX/YJG78Y4NPrBrjq20tXW1n2HdP1gSz4JveN
lsQZE0zjz/27CPx0PQuskshbeUIrJRISRi3w/Ny3E3Cikh71GQrKOGZyuQGOKmZe
lGm8mOtS324VNa38LgepidwLC7fnIm1KIUBAblcKCatpD271V1gzOQOT7Yud4t6A
FhsdlqPSu8Dp+QDcohzGH/88KatakYnhVfMKBjpmFCFUhiXsieFBpNmrV1LUJ/Vu
+/w3M1HOeNWBRdZgn/k115vlhYaOl+wbUYe0LTl4CWASBw2pmglNU6SkCgwiXuF6
RRqQxefsi4yn/CKkjIcB76K1dS0uMnrApLPHcQeTe6+TDdfCJN1SQDE2WrKGTVRI
N+EaPfflXWBd8seg7+55p4aYqujYRZExjt6eZvh/EZT7BgWJa3rTcjJUvRaMw5pK
G0SexyeHQouZ/AQQPPMs79uho8pj0dPhdcELEPuES1DHUEHllQ9OVbRNiPXhubju
a44YzZcYe356agq3K7AYkuuiTrBdCiGr0eCPSYBM9dmjg4pjoyM+KUk7M0pFdBNH
x0StmZPYqvkMxf8ZUkwPn+hQeAkuDdtTKbBb8WN0msyO9k6nud37MugJsd5oPKYU
db9ZPpZdtiRjF8VsgjFDIJ3rCNZoLbVtwzCbaDnIsiyUDH3dI/laMMQ1/mQhoyKL
jn1lWHm5v1TKVid0XJaPfb6gtJl9MfyZsbyPqZla3ynNo/ZjWCYd+6Tv1q+nQawi
D873BWiLT10whmGyFi3Ld7Lr/tz8wWERAaCYvy/epS50/HcAPFRzymOwfM7zYauM
vLLiClVZwbgK2fwIlOwmXPtMG945aNS2z8wXBQO2de6g3l0thqGu/f3J3nl1k0Tj
9ANEuQeTtVzqP93XGMiVKA==
`protect END_PROTECTED
