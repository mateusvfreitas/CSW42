`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
9YXn/dt4B/5rVUXxj3B/uptOxL3A22FTw7unvBj3iNFINiydRJpuQUvhVnjArTyU
2F4lUOsDdW30wZcC4iH2V/jugOOv1NB+kbTeOCrsj57l177/gTg5yq2ybgJAqwRQ
WDn+yJWMflnGvhwYcTrNZvGq/WhZDNBohAC79hPPzTEEMKlY8ZPp/7kOfpxSDNp5
A0r6h79kG0YNhHOH0nBvuwJPSq+O/UOlEaZsYBRyjIwIVL7EW+Mhkh4nPBFTY9Si
Q4p/CWW7focwFs76znjpO2thlsQC5aKQud1ZkO4elC9+Eu/GaCjn6EXgu+DP13u0
6dwMUaDYscomuwLFHpKxQqaI8zyS2AnlFfkT20bx7Se52OZh6510Ok3KSC/nLfeH
xdrSJvmPLZswDAnG7Z/bm3IAvirpxyJUG/R2mwawDVgI6V6MwPE0DaOhk1pdGL31
KlOkWrqPhxf1SjVMW5AAuq2nWTZcqM7NsNmi1GIl9CbE65YDrIF8hQZuDDgbzkBC
9f01y88NFyx2lRHPcvweFAudo5Wo/npqNFmq7ajfhYRpbHFpNH8VO1k8NUWO2MiN
+m69YTRpXieC8dODCUJ8uRdy/xlBXb+dIR18PDPJwIR+4ADfUpwITpd6yGlsTw9u
n1q0NcRfgAQKHzQl+yd+GOptYlekrTOfZKDZTRgXfkTIY+Vx/O19Yj0+9zJY+vtz
xzbVKTKtjMTewfbMMvfVY+BDmL/XyZPZgTKBGT2xw7Esn3OC/oKq+E/VTKw5sty+
yFQkNB2RDij2891qE4XwkHuIdW9P9o8ssUNLR2DQrJ5TVCkdEOD96nMXMBjI2vLh
pLt0Rn60AFL0AqQeLPYoO4CJqdZ7/py5VVNZBSS9GI7T3j3uCejRea6cVjOZI3yp
WU82sExIY3SS5io+/lpF3h8H5j+2ibMkOlarMVRUQQfpMazFZeth3h7wZJHBHveJ
mRyIRc4te1CnVCpnvAs6A7xqwJmnMt6GWuzlKfnp1cNiPbOOac9w63ReXz2UsQT8
UFpSNatRMiQeTf0OnS2pae7cV9tdaPlwiHWwpQd5cT31LB3NaFxeh3GNHFjE7oiL
UnvKIv0pvgyAfCrkUMef/fKQ2Mi6LYyPH3IR03Yx24weoWU4s0pJHlRXOr2L+JRk
bleluKvVmQRR0v63kV5MKeODtECDP+dhM/au/nf9Lbdc62UVMrurVQnng7etEziD
xRU2yE34Y2Wot8cUIaG/zmVrSt09cyKy1uLzI18xqOr2u2QS7gXUnbey/eB8VNQv
7AJYZl0+J9XOZ5h16ka4TrBNOTujebd+UuwNXZQTkUUljbmtwf5x2MRUo1StkISe
T7xX+M4SVWHRfhlKO/LxLrzLkzvFMlzcVnjjyz7iIEr9mH2iLoNbcQhFgq5USieb
5zwD84Sm9jkwNxoQy2ylDFQbqjhu2mjx2v+hKR4a8pTG0od9vHW0m2F+LGyFseJe
f0P+ohhlR1UFZ4FE5vy+aq57g3kOxL7906mvkNyNK9h6+bUmF8OnQfymJ7bLBWs7
k/7K/9EoGdGC5mfdYaUB/hDpUeNp8Kusbnop782NQq8Usa8cR2cN6BNDebkct5Ol
5OBDCemF2KTQu4DTOu6+Y38/b3DvS1sZfzA55QC+svaSdCuWH0CZAlQNS1W/99+u
M/ZGydD1ayARFpduo3B75Xzr5YP80rTunsg6RTEEhzztogJO8sG2cK40fXr4P+je
8umNygfvrSljyMaz/fJrrGKqHKyjmzLcR0YsQ1a2cK2h0ND7gh22mDPImYAmOB54
KNo6KGSc30r6TpF7N1CfscBuHKty+gILTbndbtyoHUaIGo6xmEKYHPz22+GXZsHZ
7U4PuUcZegxjk7eGJ9U6tegVER2B2QGkINBSU+cQMwzItyGqE5jrU+viObfQ4jvK
zIHfsEODD0kY8wVdjW/fOxEZWexSCiFPTVGqiLrkLuHdxv7dPT3k2WpRMjEyYrS9
7vrWpPH/LaoNOHfizEYOvhg9JpzeA1ks826dmn6cpo9EqKbYs1FI7JCdsUTVIZ9x
25Yr6wjz0ASgOxBXI7oYODrM3Gzzucb+GEdVO3LjQDI4E44mavZjx2KHEdPMeTey
QiSlYY0kaR+JHWuITn5Elqk+7eC1xQs6LENkwUV9cbLKP2dSCM00L6MqvWyub7Zv
dluucb3PLy0dT6bnftjw3Nw0qQ+skmPwxdk7Yc7OgPx6Z+sDWWgDj4JrsMn6Radd
4Crg6tDSw1DEFr6+3O8Z2Y53yYoivXO/3uLiuA9kBub1NHjK9QC4z3baE4Gf5rqr
vI40hHbZcZnbTfXlz6ww74NEZvn2StVv/Enz23r3Z2etzeQZQQX6dN7XDmp5lj5K
X0HKH4p7DfxcECXQZvlploZ7FfWLbrEOyT7yV+HtWmEWmVUlrbl8k3ZSiumXLrzF
uOrXh8exGv4ybkK76NdYwRUwd5x4hgfszQ/r4ngfejys8qH4xX28QI9vnWnGV/bZ
BNSl0gCCAnvOboliLkI0OYDXcvOd8Y0FNGZujCA0yMC2jUj7M254qGdX9jOH6HOp
EC68XPwFrwa7nniFCKM+KejM2o73YbBR7AWQOl3OFWbptVKVcYHNIUOr4qYM0ZXV
Z5Ck5hEiTSdr1PtEButGTJwQuX3gP7pyJYbmXQRBmN3jYCn4PLKPANk64ZvxqPzW
zbcq7/7jjJJakONDwuVw8D6L9a6dVWfLrVHXIf/vwRCEGtSghQRd7mGhHb74gCSf
SKTUZ67IyqoZj2cSLjrBwX1j4YhtipO/XaV13KZEu2skkStgAKTVLzqvu3EhGXwW
cYyqSlKHD4v12mUixL/+gOJR+UF99D3AQ/Fc6qAX2KsQeKXZ4TGa1P3vNrCFC3W1
Z5OHBL1X8RsWBbbzD7jFy8U0+G7XvwmGjlz6G36xahUu3H5QpxTz2gmlcVJrKNwt
EVInKZL9HZ86hVwHhk49kBPYsIG2FVmYn+VbEXR68zFqtGogKAt0kluxZ+Z9ik9R
nxay214TuzlD5FqgqU9+zUOezOb3Tfc8hV9PXDwRJGyCdsnv72mjdh9fgAeT1Cwa
YxYTPpWv10xGHLYfETz0nuPjQRfZFRfPtIxiGXGSNBC7Enhq4KUZ0SUCf8mejt0X
eUkMb3wtMdT2r73HG+rDwcGKtA/z6zm51D6Do8lQWL6uryPuYlZ5CbF5St/Snor7
qhWSQ/iGR/FprIbpXkqALHW3RheBerLChhrVcph9y2y2Jggjz1ozyrYB4m+En9yi
5eCY7LVx3JNbMr4vyG6a2kckO8Erhd682dc+LUUKnkWmdQ4NnqpUu2qB8visfPRH
kscVPSlvtZNMPOfvvyS/ds5fEjdPW4B98fMpcmQ92ZY/JusJT7U+HJ0E/CHhastu
uChxcVsACjYCB/ax6V7rAtdpFLk/qhTF+PptX4GwSwc4hTa+2aIhE7VmqEGNh5cK
0gZmWy9W+I5jce8SsRE1cyvEhy81RztfvrUHTDrNBRmPtxdIQS83ZkadX8xEF9Kp
CuAYmATnsa2Q7fMhMESpWINKL2oZKEz5ApxE7qzwjv1F+W4EPscWYrK+4DljCXvZ
dpRrnSK5O/ebD1WsywEnknAJoCLH2K2m1zfOkiybdyjR8zyQGx2Lm7E6EiyWWNo1
vBMPdAsRzYLWpUaF2v/9vK8wq8qGmqurJjUiHhfIq/NZG77drFnO/LrhHJ0MUaeL
eDg9fnbQAk0XdeisPHoyMHOpOE6MLJNY2bRR3I49DcyftKjMw0yMx+rOrXQGKNAq
UKLaVMzEbEqfYPN8OrISZsA8n2CHkizQJIIbwOdsY/RX93Y1bfPbk1ArUItbFdjl
MX3NBroVqLLgvMTO5kx3OeKS9qPjXmcuE4xi75hKrDGQ8JgEobVUoVE6/6PDvIaO
6XQnl6z/zN7LWP8PCSRgfNix1ilZ8b4GwtIuMSwOqB7+/3vpCXk17y2T2ifeSicN
54To8Jd4z4Iuloc0kgPP4U/p2t12XFxesgVxan3/UDJUS7lKZEfZCkauNhqFlVWw
bx2sYC4gZf7HsD2i7jkl2XEATKF5NfJi78JO7ovMXSlu6arDV/BUwlQHNf6CH8m+
Ovgr696mTSIBBD9g1CSo5rZSODM/gEAz6cVCsq6AxpZUeJ7k9igMWv461h9mH6NG
Ch/bH+EyosXZnmALGTnzzkGEz1AOVhC20hSnf3WARQC/uCc2QJuwVc0zPXYJJ+Ju
wDdj6IXTE+w4gVf+n3QwLn2POv2lub/Xbk/XrE/L+5N4qjlHtWc6f3F3U6A9ZJZV
vlsQLXo/yBjoeViEfB5fMhXnbR03NLI7l4vsK0zE45wV2OQn5rjoZme/0w3AjwPB
QNk7s+iMCQk/AvMQoEBPhvIyRsI1lHmlhjK682hr4cSISOJawBufzPiy098YWy9g
JSSWWk43buAsNShKsJ3xyD77FIWAsJgW/Ci1tzye0K9Ca9BK/9PyLuFquR6JIn7y
e7n7KP38i8s8DcECfq8cvzbXrCs9TA3MPnO9zF5KSilpfflg3nKQe8S61TVjdi0C
ZpFAojsw7mDAnmKjWKenxRoeQIWU0efXd4UdW/iPkX+OEofeg5WlzvXcrrQLKC5A
rc9GqZrXJ3/7/vvqJGesRPKQUkDQWvCYwaCHQ/EBFyE7UUMSiOb3Bmu9Ts595+qc
S5lh9coxfp1zLb1eJgHtKeWS767A3ydf72A43bLpbwsP3dZ1p7buThexRsK4Ov77
Q5bLVOp1o7OMaJqyY3uCobCPscVwBXfOp/BP4Mp/Jdb/1G2HbGLGVEzBPp4Y4UY+
acaPsDMjSUWKygm51zvBKaFnC9IqM+8C6oFOuzCvLFcAd0v54bh5hTLkhyXiw0WS
UxXJQbiCW2i3/JvMgY0eULOAJa2s9XS3CUCtyh8gt9RD+w001LESHPQLibOUugvE
QYHisXbWSq/vZ0bDZanWqtgbZGYajLxJ/e6SBskMGZlqOGY0gFG1/ZAZGrvJEhyU
uD9wnMEa89+EEVcbM/DnC8jP1K5v1L4KE3tfDIhwzoJxVEDuojSU5fwpIZTnatOo
pyJJGRgq8uYcBI44FNxnE/f108LkIv0fAQQhGvMlbTKsBa/VlRoV8S2DSjclusmm
2iN43ZfGG/wWynVy25TpeElE8QB1SbYPKctq+shVJVgXRcZ7zNlOHwAj6kbqqich
Gv0xj9GAg5LVtSvkfw84fljIeG0NgY52qgfAyJfJ3BLhGbrLWER6yWl5dCLqUj6g
F+YKu8cxWEiNHuBCNNgLs7vFx6QS9g9RD7ngwDTPSVSTecJbBMjBK/v342VDnxT4
LFZicMQMulU6W9mtXh2IZVm+3VYZPm5zMbSQYg9SOjmO59o2i9Mhp02itfcQL5f/
SQuHmGMOvjHPaGhxBAASaflTF4D0e2hpbp4bUPQgA0vyRAWlAgR9+suC4NRV51wx
LqQAO+BDM1LmfnR5xv73IiZIdHw6u7DnbuTX/LUh/vr/X1VYIcjuxOFGKhLpkiCX
pVloy9krJjx9sLFEGCD395iLkEti0sTpTSY2klev9w1/n6PKPrSfC+GSpKuS/+7O
J0xaox7N6VZyo8aQJoOrBXXPWX25l1OwpAw2xDrs3r6zJEZZMdeWpF3cvpbrGSxP
HoLiGzbECgK2SZKYMXuaSebqhbM9FsGLX8/Ue8YkOgiae7dOju+Uvk95HZc/ZQNQ
XCwzVpioTrxeZWjH9diOdS3wK8uKaXeTl+cILR5sWUW3ydAvD3am6AJRmobEzn/G
85a3OyMp1VS6MUC7VOdJW8R3lHnKEaJGnPN3o5qW+afHvth7odIVPqGlTm5NvhYr
0WJtEsol4N1iiq3l3WKJUw++WPg4iacUk5Wd5qAZsM7a+IQzN2np/KZ2FJW4wAXf
dzHRr3/O69/eA06ViLdJpBPqVt9b2b87y4kfqI7XY82Hg50gW+eQ37qSu7F9kO3L
iKmxlouR9Sg62lH3+T+StiMD3ngf1igkSnl14VexUaXRx/9fXx+mTvqElzZKEUn/
TcLgbGmOncaT91qQ39TJcHjOpLfBHS3fMOFjZ4wXMESGSZ9cA3nTMAZFzU0lh9gd
TrSDyltH5WRvJtI1dCbTqXC76i9zNrp+Ja9JnXrDjGGO2k0s+oos3247C2H4GW1D
ITE0ibmOFvf0jp3k5A5gfN42kTYQXW8oP1I7MgTmPomzM3NVuthkZT4VZNqG7V9C
nlPF5+SeC8D8yZcep9hwapJx7QsUgKKO1akZm1wjEk8yuDtTDDuhQ9DfvYcyocuD
f5STF8rLIHJ97X564dTd44Udck3v9n5HyjukrLuB2sm6m20NEcROuXb/LRqyhM4p
iqjUAd78ebWyjJTHJps31/rcFVXmakiUV3FLo/T1jrDR7xxCoomyLvrJNvKHybt4
MqQ6OBK1z7ZI7L1CXE8Y+W6DNRyxhoI6kfUbxDV1T5ggnXsAmcllfSJg5puSArWH
JgQ2uSj7QlBkkeQ6hfbFMFgFidDMS5HpqPy7SsCQBb8Tfxiz7pQMKmY6zAjztswE
2PfPzL/uCU0tsIoQkrwq36LvAE5BVGr5EKi081MjSCUpzD/VYu/h/bYpFz+C36/t
YZzgLzkYKS/RtjnMlYIY5ONSZwvZ3nVQiWiy5Cg++F0lPen89GOp2qDMnXJU3Dyc
Q3bFTeZutiBuk3l3qb7NPosAQjSbNYTHR16ZRFRZFyk=
`protect END_PROTECTED
