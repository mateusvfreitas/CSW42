`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ixin7cmsEvabhhhyBQeSX4InUB7Epp2gMuwtZQexOMwoVrktl8U/0Pc/AKyuYq/F
TeqyrDvaWsmtrEHnOKjyOth0GgC2c07RWGk9Dig78gkTxCV1H4Pw98i81AnykSWG
brLgKNREJV4mkAb97RcrqzMxtIy4NmBpzyKMqvZmls36D76Kkve9XSmvBJ56gLrB
EfNb62ASMuuEcpavdnNx0p+yB2+A7Yvh6YTT9CdOC15g2ce5Xe2hC4GxW0rA7bnV
Gg8oc1Ou1QjHEfLts5zoJTCg6l4yOujUpXrxLZ9rZAnyYXL1/bZ/3CbxYjki+Q6T
ZQA10bGiIJ3m7m2b/CT0wJE0QuCh5l0gTxSFalC/DDhj9wmlpOz/WJbW8VWwVJMC
5wG8F+MaSLA9pD9FOhfDfxCvY7xP0+9NN6wssSzgTToth5TuFx6QLKyKUWIv/Mxf
88LXekEx54ib0gei7XlNN+yDTi4cY6ReJOkEk6YomBtFutyJ/Ys8k9AgiR1BwnQV
X/j7KZf3gMLL58/Z/CS+oa43cctLVRsxloBBlQwDssRe5UpSb2UAwHYYPT9OHfEj
XIR2YsMR/OTQvAEP7PJflq3Yhxn67e/iLTRjUPtToOsdv0Yxs5es5lbPSVrqK1oo
iW9Ol9l1niBW8nCyMrfvSVFMQq8k42tpt4+2zYAoN80WheulD1JtqManyF2i+n6O
i4A6WU94+8+Ri5IJcOyDDM/fgkih/bDV47vDwX8si8C/9i+5kwbJ8KCcFS4ggJXS
GufHtBbDAVr6w/mMLLxijc1SQ9xPN/NkAuCBSraqIDcDz49J0SdmxTjmRdMjLpTg
5hIgjMfgbgvl3Cb+GNb/UmnYaQKvKScpRBRoM9r2znJvx0SAhe9PIqQ1mY9vR8xp
jf07lVXzs+ujYCtqiueMthVPrlOlhLOyQCGRXU0b44ReLhkTu8VeJ4bAgwEliZWT
69tCctGN5L+bCagn1dKgz4jCvSPrSjjxIsROEH6qyWs7y5Dw0hhn76IWtAhtp8hY
sMz4Ae5GcaxPEaNYmYdWzgfofAPFVExG1ukfpj1DcNPuIQXxWtnxNDZaaXqFIW7F
No1wDT9luLFwCHebCACCw+4ESzVorVNJjcysH3hLggPlVGZN4/0wN4aX5cOvtiq5
YPyHNstK1RPxzTC43vVavdWLf7sAWI4N56UlOPXWAREUt16BJd4yQe2SJC/pw0VB
RCqr8Yg4r+skaWwLdD5d5wYgg5sMaDAjbvtV2Ya+6hOgyfv2R2YpGtG/6DxBpPx0
RaGErcIpS7zhLzMU1SVeVNdq8JSYfMtZXNPhfa5gPzmYl/U01gmZ+EOL0wYSJTkP
ywhvGauVO7BZJ0sA25eAmJVI2kYyRA7ONWIHCJPIxBKQLeng5R0jDdIFcO06CNja
qBJzCesK1j3poEH7/uNpddhXmo5JF76AXsskrS2jya9WJVAr5tOcyIbaIXhv9FAm
lq7l3FcYkiDNXmLlUVxeUn0q5Tn0xTwDdbIYKJG5IjThOlTVbGRF5YLrg6wM3hNV
hHp4t54oCeeIP352rh3hPngNqKimroVJZeRNoGVFx8kLpbUfR2xw0M4T+CVS6p3m
p8uBKD+sXNbpobnNmKVNtojmxHokXlLSh5AAHjbbKumKQD7AjkC/iNmYV+9W8XNW
BGhUkhDjaaOp4tKLJCxhdYvUrO5COhw1JY1JeAWE5xGILp4b2Q3ly9/NFeM/8ISC
P3NJywPxOyDQnOpTcBqaM85hh9X6t3MVakYq1sdVPg8ok4SdFq8cKz3w4uvjGUV4
yJhwjJYyvGQtjz1PDq1fD/arvSQ5qnRjPTn1X7UvGCwca8UtaBag9Vh2L4gZUdHS
k7FcggERyxokoaVCm/lkRmoEV1zwxO08qPBlb7WR+tUGA0ZnkOp9I5f91yC4LuRz
X30Jj7QC94ad0Q2QJLY0hWiuVzqctQFHjWxeDrmVTMqdbzyBhpEpR2isrLocFFfX
um/3+nv4U3eZa/PVDOg2XZN+y30AardfwIa886d/VwKA+85MLcAEqenpR0GwS5yk
zvzRdlkYu0zWfw7ZibQWpNwsdOdhQXjY6tg1BArYEg6IliRYIBt6AH6Hl84ppBHn
TeKpg+u9SY/79fizxk+6XugDQYWpPY1yWDle/kF5choG8vSMaQNcShaPariLyfoy
RLR1k+WBsW+R1E6ZaIwpHKdBDIsCqQDZwUZ7bH5tJJ0rLqQyEWIo0XCNkOqoIpUX
m7QD+tZbiqBefom2Y8EnvIb0yBIpfjm3RNaMTTmBCmRg16RsWYWEobiojL5u3T4y
wgvO9HLGiaTqWTHr9v5oUeIYIj4wTmHb9oM7lY37+ngZHsx9NvZF5H+H0PHP+5e7
ow/yomac5ZkQlf1bvBtI78haL8oGjCXTanSDb5oY3ylopEiuhnsyIal/ZN8n94iU
Is5B2dEVWP+DCQYdoAP7934VCTSwUa76cAe17X2KGjeCsGgI5c8V0EzgG5y7Sx+p
Bg8ugzJgd8Cc89a5cCgnl1hjCaGKFICTM9SJgxNb2ZtIZAwOLnx+W5v0375zoh0n
v9mvwgoEDbvKMqCqXup1Jek9wyptdi0FdwReY9O1mP7G9ndFMu61zVsdozMbTHu2
Oc2v8Mh+PvFs5n9VK/JpKU93PaCtUMGsfJYlOQCFbqo8Pq/dRdZJ1KimhWg2XYUn
XP6e5B7Kh5avr9mb+V8I6jXNdRLxG4hdQk04HOFp3Nwuz2AKcweNBhqwlPGxvPgX
dlpYR7YQeeDYSkwLXBTbaQyCFeEyXh/Pvi0YC92wLfKlsyzms3KnqgOyDJtEStD9
wovsuJJh/TOXt7tinSHe5jE2WU/PbDVMkaqjxXZHBaNQdKRzUm5cfT4Ybf2RnA7h
/SNZ1LuI5F1Qo1e6WGgTs1iKXpuVI8884xghm4FAjgu7qUGTnW8CGrRB4vDy3b9M
odkprpEUSBf/567okB4M8gYi/iBmEJABQwoL3YoYlI7K1oIcZdIkYm8+6dsD8aHW
MQAsyU2xZgcDVyg8rwLI8Pilede32WjwKznYr2iYOKCqtGRkLSUyp+Ym4xQBbjuA
J2AmZzrIaBDT5cjbilaFuqFtPiuyUx/Yr0mhqkklDOvk17VPZTWO8BkuI7dIpuuh
C9zwOcBaS6hp8I/0k9REKpsZKxOI5cKMjNIVwcGVPQd+qc32c4sUhR3GwP9Ry12A
+m9AggRkWrSfaQJywIY/7wM8uPoPBtA0AwP/OLe7HdVJO7LvloMVpElNKqmSSasl
HU5RhBpwRlLbU69C2XEDa6yPx7g9A3s6ru/e5dQSp/LIzZy6EHlR6nCEs88HRYJe
25aT2VPYaVs19mJF0buK/sOgg8lOdbYzUdb87hiB0gJJJoS+kXXb5stYBVDxfdDL
ekOTo1BoPQxU+AbrPLT1iSjuvw5zl52SjD5vsdPPl6CIS6OlimQ25BYIflLOFdgV
FVvGeVJuup284TvM354FrcE2zh6PwFKxMhPIWptuRvwDQvvJBsrNkeE3V8nXg/K/
qMWguMqPlvqI5ijLC8CuCIA6YbrhSdeHd4jWD1N8sm1G/TiQ2Jb54Kup3EMO7Hhr
+N81LsYlyxJsQ5J7gCMjSLddF4JOc5uXZ8aTzwBMIBGqX6d5/FJgy/35LBZd5mPT
HdlkjT+VpRPks62J6Ygo0ZIxQb4dv6hXxhBqD2WQuCDFemRnw4D353cMLH9NgNQ3
DHol3T+BzVSYyquiJdOymVirANHJ4swoNzLZ/dIpUMSYmb6iyatJvKtcLZC/9Gf3
q+MLyBMddBOfroFb4rXErRKbsZ2xWZOPyzI4Bk+FLY9YkxwakTchy0YfVLhC68d4
RPMc3tJgfBCxhXKr+2P8qg6KCvRVTr6gQIbbadnzTfJR2drOuqYhVR/lUr/+KnOs
bV+uf3umwqoSx27s6BevgF359/yGwPyyjtYy6reOyykd74MIqQsYtt/lx2FvMZMF
4BsGt6bg9FA62XbU8A2fuooOraxULxzKiTpunxfExF2J0huuj/+jsSRynGO2FWfj
DXqBATWliOPLEPCYW9PgN+qFeHex8vlMp9a1iLE2WFLTdjPSvKH3gWNvNnrX5xmw
v9avZcwAm4P6yQaHPIncahvwnF9b8cx+/cAp3ax7KzEaL24/3IoT4GfEp3qhkzxq
UL++QtgIJfMrwM0abMhGL5BCkj18dF8/Tu6xkB7tjUriXXsVUxP4LrUiBbm3gA2l
G6yVdpgu56IK3YKpKM3xsLp8dSPeh9uu2Z/wGf8tOvCUpm8qnIj0e0h4CdHyupZU
Zpg5BcpEMoFiq4o2SeiWZnRZbKDkcoomOfW2q9RJcjFkiBsNhIFgIYcrLLB0L2wD
a1EOYQy9clfOFPdpvdH7FHkhXPM0yfnfjQnAygiF6UlY0PXalM0E1Z2NC2CVxINE
/A77IUWU3rJkFBVaJw4umUYLaN71uwslREO3Ua2OKwBFCv253oatYW9EGcRHp+d8
1zF7xGj3TWI2BPu32r997Dppgvkh6hxxHMEUVgEc3jw0ODmwI4yOHt1YNjpprrCv
032rnRPa1QU4Ki86VhRvP1sYxX7hIXypY9kDxLk3tmFIqWNeKdVhrYtKazfaexUF
M4wST344bGYipyGXQ0Rhx2TuwiGqqAGawKNxDeoW78SWZt1kgk26cFxdRM2IlbSu
8cnNLW7L+TS7doFK3pkTDyExwXTkRe7knGCge2y/Y/DcflweS5rA0V2OZWnYjKKY
+9REpffg/f5sTYEBKtRv8+gh5yiwZ4K44/kXGqVq9n/+AEPr/Dcv3wP1lhBPcwz6
vCxs+jgb3r7G37Ns97VWboblaD6FDMfjwvaRGz9yXNJV30e8EcI0ITe9WrFHTgkH
o5GgDCp+hXVuBx+T+W+RE/9SyhLJS8gBrtoatqHhJJpkAm6m6zoRAWdSrobi58Ai
uEqYRlH3nNQNLnATXXIuklOt+IwVeaWaVIdnyf1LLJ7jG/tnCyo+DmbBktdx8WKz
aFY0f233wFQP1tlrsMrEQz/tboYP0MKGKlXbD1OMlW1xgZNIE1iP4aWtG6Vb8sW+
jswC0+DVzKas1qM6htC70UaWQHl2nDh8YesWzgSSMg2sq+efpI+6XxJE1D0kRkTV
TvdYL1Gbl9G4ZZWl6mD46qBhAgEC3M7ni4xhXhP1AM5FPEJLNRz+G5X8aQZOAxEH
mNy445r8QUe1BtzzylLVZJBKojlhGbtQhj/gspOmOMohBnDVLfzKNrjSd7DUZa9n
JAe1a7OO1b01EKQBQtbRkciBL0PrBjBlyvf9R8j9ssn+KGLrq3N9RgJ1fQs8+/Fu
C/nTKq2ol8lxuOudr+eIM5icvRbxAI3SDc2GqJGGF+PMFW5RE6t2U+1ktwyVyG5c
Arc7my3aVCLDkCGy+ZOvydZheeEAJRGjGIYMKZFvH81UKxJCjt3tqriJvQE3l69Z
X4hXE5DvaYgPRoAh+Tj1rumfytpDhoEOerR6YE7RvM1sct3LYELOjUyC24dPvnc8
Wl+Qd4DUTNIwO20Ex+4ohQKeBtstWbKj2fTjz+UkVhu2gxJ4QkRQh805NzO/zm+A
Q4YciSmQpwHvXltVsR4y9ZM9Wzrgq8bPkPVKjT5qElui5NtBmTW+w9VP1jaBVe7o
ZMlMaAwoCXw6DCZzMBVRElXvDwJMc9eIXM5o/8s9wuiRDdFJAp+7gS+QwDkm3yu4
zhLnkSsTJuHkbp/sd6MmRwP1rp7XeoaGHdFHC6/myyjkYoH5B2IwEXtdaIsnr9rN
QcnghD994LK3OC5wSehO/TkeQTA5+q7nst5HcaDrsRgBPdlfOue+1LGUvqCCf7JZ
JTzBn6ZFT5mDDP0SKZk9jAzOIMaGbFDDq5B05szXiEBG+Hem6VTYQdvvlvvaplI8
469wjGki50FbeO4x9vyByAj1R9caM1THrH8+CwcswEHQneShSFZFv9OYSNISyYUA
i0Th+5JYWAHPqpVMrc5aGnr99iLOCtBMF0dYbvizUfXIAnkvyXcK8RV5QiXxwnpn
6VWwXwOfohaR4/A0phzrDvGxmmmSyVkKaDd8sPh112+6TzUHrWsGTOzusV77VbfU
axTK3nxEIkNNIFwSWwx9lRougkifXdHKFGfOQHQfKp8o2/1f0qD+Rp6dRtoNIsfc
Uz6ArpZ2aFd8X5HQ9W+t8BT65zPUUtKkdgq7fc4mpMJ++KsqvmbP+QSCsLFSZ3OO
tYgP8Va/q7CJyBdSxyD9ZOpHMdwx+p58UH1y7eUQFeJR//Z+LfgtaeqdRDmwyGER
y13BtzXNBwqDhRtMi4UCSt3ASKEpP28mx38etHKtZvmH9oK74N1nauJL4G6zRGQ2
NY1gGEhsVcuPChVezJU9S0izaOSeUjZWlSEzDEq569ixcUF9OZV6Bx/Ub/NBvBbN
zTQV3Dnx9UZ3l72p/LSxn6SzKbV2vZIZHHpixOO1ODpLkOHYRtGdMl8IQhE60w2U
qIBH+iZyYbEG1SfPsHPgAeQZtw6jo5LIfdOJ/8qOUvEy0OQEWaM1kmlMpf+RKr5x
vlJFcZw41tqgsdWAWCOrCYAmGVN2AMZn2LALVGHje0rdTC6jpVjOAZqfzbRTjIhY
sQz7zVZCDplbUaYbaw/Qjj16cqUp0G5+7QjiMDNFBovxLWFNkE46sa6c4p5zUiFy
v/tbomuA8dj8cUM9VSyZs2inTGsQbvXLbTwEUO4g594Cb6OUFs0lneot7f0f8HNd
LERxFKgNchXOJttY1XbS5OHZ+SaDCOCl3Tvo8XMMfnCg+biz2FnA70PUjf1CFlaK
RcRJCVIf54CbAqJ4mqRbc3L9XQyzrdFJS2B8tR+TBD1yL7zC9fXn21sY8Fjp9HVZ
8HzBkT+pVuyfWyv/N7bV2ONkiLld9cQimZqA+JqvXa+cYvoxMDYzVAfu1PxkqRri
odLcA5CdOf9OLHkXeO55GXYur0H8ODtu2zJryupo7EOJlkDeHBg2XbBKrqUHWy6Q
XqRibsDccuoH7v/qCDArBVlECReh0BXT+5gpQVZyZAdAt++lbgSpzxdd20l9BcJo
XTU1XlgkJ77z1K4JvDslBNA7JHC6UrX277wxXQ5XPFVY8VjnAuFQjhURnKnSf/07
YwdSJCyy4yEJllE0E/i33olZRnTycpiIBDne55MmmMv+N+0CSeMnYet4ORDc1aAw
5BihHp/BXj4pw7hvD9RhAaPdUJLp1s+pcqFrAVnDPKGRSuQuYrGbs03plVyxCnfw
aIwdMrsyXNFfqYT3hS36WoBR3eoFu4yLFLykU4TW4Jl9wVReFJreRq+Q46/guO6z
v3IFvDgl8BzXiMIfuKb8B1kVP/D59j7LGf8MR/ApjALhDoVdIiaPF3gtSGhK9VTp
EPiQ9WaBaz+MvRG1SGHqe7WHF7krAfHf8XWurS2hbgX8M2UK1dyCeqSNqilG4YVT
UhuBml5nDLqy6lR3VS5d5Gz+WBbAb6/4w46RMP1UFAJM8UIpdjOwPz52gGbWml86
bojUMVr/mF7ghX2IO25vXftDYOzkTtZ/1ioMwnLBBixiACnW831wJs4DsjDOY3GA
a00mJufLAz1WsSZUbgh/r+95SV2JbcD4ZEfOfDkeYjOu6yKBy+RrnkT7WBPaeblq
dsfsLMsEBNy8S/UCTFPofbGA9o0FeylEx/H8zuxIQdiee+2MqsPEF9MXuj31nMC7
h1p2w9C/5afo0dFuMGMhzCpaw+HAgGNJpjxbvWyBwssbOM+SMQcV906ZSDF9lFkI
nI8agzZY/LW8Sx0wMbdnyeZj4AStdz+8q0MYhw98gQ8AdRBkGl6t7vFbdB/wO7Ur
4RbbY1zeDVTKqLMP69ZyYmG+b0uDsW/92/H3JaK1zmrqj5olPhGeFmtsd7dnWVtq
jzS1GHh6+qD/Z3mYhEDb63P79A8BUHtwCQaWrTh6a+c+RHXuhgc4e6TPumHbO8S+
7iJI3qy6bgu23Ep8eO2Y0mRMP3BmRhGslcZrVIiIXbNvDoNwH5iSRptyvFMIOW4t
R3u2J7cHwRRSKxjQe3La0taNCfWYhoJfpAG57ywnrYbUF+i3qECY8TiadCzCXAzv
jZj6zsLidiy3QNF/WvE4fYNN0l5Z/jIGZy59QBi705Ak04Oa7CF1CzwIHxh+dTsu
YH7C1N2jYiZ8PhFt4wR0ysV7aboCFM1Qk1AqKfVwoS15hlkJb9OmnY3Lq97c7Dyb
vZCyQIqpFGC/qHqdQKhC5T176iJH6TiQBimGUQc9OKuzvUUFCYapG5beGQq+iCZx
4Xjmq5vgnxhcfuDluHe+3zFhwi43oUoTzPE+DJCAHgW6hYc34Tne673C5ixRb1/E
7q0e2Xkrh7fGUfQKe2636EBpOudaGgZHMfJFDG/rFglHennbFgqrci0JJm7nTEQK
+Q28xDmmS4/0tyOfYt775mpSzFKCsePZEqFIehLV4nRM2f8qvg80li+l9WLXeIkL
GlQDhiSndNWoaErxur4NvKvVfHAhCGJRIPjz/XY0H8I5Q+2ekEjIesRzOdR1YmWM
8MqmpRet55ZgDIKxKXCUIZ7mzq1nQQeLn0BqqcagDK9POKhldxRolM5E25+nPSOe
RhX8nlHnbTd9ja7DY79FCSEbRSeKsgd4ePZjX1OJ5h+CmnODQJ3CbV/C6TME3wMK
kIpYnNGOUC7Fi/4IYqpoF5SdCd3tH62rmcNJ5u62XH3h9dMAeRfjToRi0xFosCpx
13Zt6asA8XaOm+5MIASp38/O45VBVjT89bY3Fu+78LhsdF1bQBmPNUYxu6c78kn7
2cJhrjdP4Zw7CIqniHKE0n/AxfOnyWTiEUGzpHeKz9PM8sfIJXPgT924ekduFIiQ
IYMqsT/Y9VzsDWCSXeY2s1a44GXm3l0klgo4H7sewi8JsMFJ44sYxidzbpqS0y7k
JkyUEaD+8AMeaDQEJTBpkYac2GJF5tChSFebqge4rhkULBX0v1vzAkhY3xlY4Hmh
oM2uf2CmPzl/DvmA22n2udqnZDqKzqu/97YEKNRoKmyH+LGhpHg2Znn4b0dzXXxr
VLO2ERHVL/CUU7TiSwIlWtdBaCBD96wWFpEE+2i+p0U05jfH0lwRP2xv8c7Gp/M7
ODeJAPTLfInSeaF7WyrWx3zKyedscmPjT/YVcYWKW6y15WSysiAsDzBvXl62BcKq
uBjbkVI+RoPHR8aKHRYYkh0ws1aY66vQZ9XqsBKHEthR7zVewit/acBGgMsy44ps
iV8GF+OGC6+8kewOe1GsR93jZTFeBir1HsWqhRgKxnIjA+c3vKsUH7wui3ud+Epb
G26UUTiKlMTcfMCZI4LY2Di5qQVyeRZzD07120tN2CCeNWLlK8NDrRmw4CoGRAu/
0oTK1Vzj7GxqTfF3slTIKbyV+QxT04/Asq0MRco4xmi2uZ4XRWHTuMA/BfQYjr+Q
7eTD7u+Qk2SJzKxttevyw+KD1jz512K6RuZnFXcbU0kSbUYaLrHG3G+Skj9nlPaO
UEfbrQTqB384jjgkA+Pf7LM07f3XoYwP9MeRhfhvb8duibSTPVGLqO4EORry7gRQ
mzWc+GWHY0a9mpOUa3ev0xPQKVah2DtHIaG63cNRQ85fnXygR7lrPcLPB6DxvsZi
EWXVI3/O2I9LIru9WdllBReuNxI95rC0v9Xi8TTlbmdSNuBodTkjklHFVIzCmwCF
9dzrto7LICO5XMIgn9d87SRNIDLUmi28p40B73/pgHruGEwBSo+OFMXsHjXJ61Sm
JEJ80pnMNOGybeOBxncVUPH4v2FI/HWwxxNoxkzlQB5fLn61Bd3YLx69TGEk0bRO
CMeaGCs71wSvMhqlwovpqqT0w5YczhzzX0mOrkkEnEl5EA7DYgccI0YLCsgnhgqI
8Q8H0uJPNji/jxOiYK/6Z7sgS9V/XbwEIk2In4VUBX8Niswy8OTdOhIqkddmN+z+
RoQxGvfyXu/8RoxnMy8mQbYgW3tyvy3MKHI2hnZCAtsCiuOfi7Mp4dHkDEdryWGl
ILU14cbYeJHUSZOT7OTAnpO6/3ykME8NB9rW6VohG9/srTrmH5I5ZBIEY+TnxAyc
3QwAeqvFa1yNY8sqSakp/Cr5RQBWnOU/OplwJyZlTKyA2m4E6Z1Hkcfq6T+VUOTi
kepnvFHSIUtCuwBZEGFCWsNcWcjHTT6D5OqxZUlitEkRqXDLBeZiqxt5VkCDm0P3
lVFAmX3Vp2PK/l9kzrtryo9otst5f5VyUkLwvdcNV+BiokCS+fbPHmr3uaeXSRbA
qrYQBGp6hGkeNsiEOJ2pZ5ZJ+/Frihg/bZkd5rk9t9gUYo9hT0sLnvWY4mIWlI7Q
TkHBEQoerq+bB/XNFcPcpGJJNvQBrupPGhQHAxT8BlwbytLssZ2j++pNSO9WwVVm
DW49kczHW/3Z37tMaMWF5jjCNWdmfJiMAlGkzoPy0A5FVSPjXcPRGJNPs0CxYcq1
3PRuXQmtBr1xseeSRW0TaBaf0hB3Zw3I3Eu8yFUbgpc=
`protect END_PROTECTED
