`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hCSkmaFTMtC3l6dNqQBLhdzgGf8DlbdgUraE09Xdt4xBP3XmY9EpOeDyGh0VJ3gP
wgAPrlO8sTalDvT0Vqhrq6Eyf8QU2rG2JCXRbhi2V/WJk2YRuIhVxV+o9P4Hi2Gk
yuSgLwsG5SqzFPthAEfGRpLR8moQjtNM6RZEWc7FYVydAhScvjEEyklsx8S/AVBK
+I1jxWKaGm1hVBTgVnetbxbOG03cX8gYl3gF9Tel3FeqmpJs+qwVSri+/95l18xZ
nOtSLc+W5x9RW1WpPH2E7GLlJRQopuCeqBFO0wDpLbof4iDRc4Y7N2XxoPBRsh7M
vmSTNil5ySkPCKtzBVOxUBoj5wovMz/XQllJpL+Izc43g/immQvG7Ur7QzrfF5mw
Wko6d7E8NaBOJbtj07PzlHVEj3MkTCMrDUnJu5Rk0b3GfWSlPKsK3OAEzEuPZ1TT
2aPsxsR3rD9obdRr3gTH/k9597DYptsuZKJM4BN0jLu7/DMtjoNpxz3CdgqWe0Mi
eLrxITa7zztK9hF8i9XtNgwE/f2XiMveGvlhoJn1e+teqnNnMFCmcdUfdw330fXo
G/DkBsAonwhJmf400XQFY65lOE8KD+cA/LBXfFeEVE6DBajvzkbPnaAGaGSO8FIl
g4mrPgH9a9jQLVi1RU5gCY+TBFDp1UVG5e46QgJCwHxdEv/X9Z4GoSePWmdk6nD2
fJHJIKRuVgRJ6vbkxPjTGgQkNUpA35AorPNIoPFoL92f99IBmp4BPqvewPJy1/Ik
YstuNadiYhkjG6hp3AJrCJMJXBjVhyEjCRof+uDzWfJ9n9mRNTDv6+938rTi6/bp
muPRlMSOyOav1AefX1WoaqwofADalzU7Lgq32Fs3hxg8MHNXNAClr5IlClIoTdEs
YOpY5bOhuDk/BSfnubDfk9t4+4gQ0rC5zTwZ3cuFrZYUyhcEGlGuQabglViwIDdQ
xQy5g0Rfn5Q3m8vPRlVnVQq2ijDavAAa1K/7a1NAfOz8fxI9CHQoWjAnXM5JXHJW
cNePvsJTwzE6Tbxg4SGNsWB+j9IGUbNoYT84vRDY/RX7XciiDCTanStEGMTn7CDE
ctfKVJLGAcBCopDr+Jrt7OuPWnXwF3+TwtWYR9p/lUHXqxvnS8nulOLWcxM8fIyd
3ssauTVKEF3jgO22+78GJWEyb9N8QIrbIZ38ETWC/cyVrPTPCccqWJ5GbC2+lhSa
COdM/Lx2OOwYrlR8mqj6tlEqS6U4kOlfAVtxN1kPAi/GtexqH0YbWU5rlxA6Cp2j
s21VlUc4AT5ipjVH7wewpXskZYpe9mRLkm7QpPwfGW84oa3M+FyghQt1cJcEraOi
sKSMF1qkUaXSW7ULeGh9bJEuXlAXlRfk0n/qgIpxRcGoTPVR94UW4k9AfDST9D+S
AN5eWV0dL9dBSjP5GBAxhNG/u4osVIzuuybodhuQiK9ycVW1SEELIh35b7FRCnDY
DT7+tPY/kVV/87eY4QxbQ7jSWxf8uZJ4OzhiM0WLWrf/B119ffuJrkfvxwbnF346
D/Z8EuE2tFVkoTQHG9JOQfcoGuD1+3pn63hmkXpAZo2+sLw2KwzN6H/lw4u4DJ/x
2ZPzrbimnwb+cKqQevYj6pTU3HyRVQE5gCvrmUNNvgz5W7RYZ7PayYAhGDdA1QD6
SGHdRsfx1OArN/nDxFU35a2MZqE70MIQWf2JHg9/vXcpSD1kPn/UkRBgAdInsrGH
jQmBe3UpxHZfqjKGm2/ENQQjQvXgQ9yykMd9Oampay/MbXHmoTU+2QMxA4+8QHSC
Q69T43D9QuwloyuqiX8vyQi4UFcvyWoQp7qeYGjipb/YOr1iVgTMn2xlqcZjoS9+
FP2eUtKxmM9PUMDpqGg4oUOMoNpa0U5eseg+0HcefV3gE0zaJV2oRQD6ew4h1gbs
emjV9KY5PpjQ3WmU2WQCEXKTs7JeDJkr0Io13I8+WjSBPOXcz8JZH/ZB6UUKWzr/
W9DVbII13C3GauyCqQgrJkSbf8Jhk6/j12XoivlUWqs+9oy+E5cQ1BzyJUIwASvb
vtp1epwPrQcQwyJqFahUDYsTfwmuxWAwG4GQRzDLApcc18c9/unfIWss9tCpZ/ub
O4bkDxpv/0hiWH2ClV9nkIF/TysrfvrZEZX13qWLSnAEoLE4qCf/xeEQNykUlnLM
X4skiYimr8dZWl+aULMki4xIbFDVjE4SmyNGTW7569VtzpqgAvBzZec1vURB7pHP
WVRRv/f/SDYHvn0gKQBtQ145WICQYGEDRZJOU6o03tc23YWl0vmbQx+Jntqakwgb
t2HrZRomkujD/aIS8UUMHlHWUZeJ0oF8TIa9DR446NQ/+z2hRD9q3NtJfmynDpTv
RL7K982rXPuVyQSTxvBpkzQdoyJN4Xq2uJAMbMQcRbmre/N+G6gDRX0KLxZjLsnZ
Wvu+h+39A9f1mXUexhrtJ0IBc5G4U9dj/TzVKsySSfa/VetzAyq/q5y2lb6do5Jl
CKKCrKOy/bwMjNU2tl//JWc03bojS8ntSm+Hxeq3ESaIJNZVwKgNGTcdMXGnWglr
grPfjr8IIEwxouZ4/rKYPLe1goHw3BSp0VWB0tEFbCanq6malMxOV67nUCq9i9Vk
/xYuAUvl5Suh5Myx/e1/YQj/UApBRPTi1bgNsRtypbqiFeejmR4D9Uo7NWmmesVh
z6TBTPZuRrDGUrmTvpFnuUEzbi/+sXmcvam9TobWhDD2X6N7rec5EfwMwvNpkCXi
7ABu6U4+MKc+dI/VpVvLwDJ3Tx+Cb1ctmXX3iRHIL2AP+ad8Q4AEFIIwBv6vNZZr
qipQ7tvzm2fQzskLeXTUWE5VMJBTAEPMzkYINvi12hGShNi26qt09PQlStsy1ELm
gmzJWSblWl5JgdbsCY3x4xZrcAUsimrpf0+oxaAHmu+i0reJxnTiy8jyTCr1NXQ2
Z6Z469JrsXeSQS9XkGT4sY8ZQvzb0XxQ/Rvpx9W7/Hs5IYlMfkV0YW23CgWGADTK
z/SS8il3nNr87rmCCn3AWYtv3bW1Z0AaU69HHR6HJEnrJdSkDBrd1FAJ+f115PfH
1kbDEh8uKXW4zs5ADYmmHn/tXvnbYSowS2ztMEvGIboZjP8BuFfqHplmM68wz+28
VAqzqxUC9BeR4m3lS5ucAfp9Jdso5Q8Zhutqe7qXu3LhBcrt8s/GViOyeNZcVG8x
eY6FROYK63G1L/vu0/yaccE8r4yyGvzrdrHrWT7mIQKuv+lXcyy9rvSIRJfvPfSz
inngW2kTXjalbEtcvqavukjCNwREex3NgUh5WUrCWCnMltPcQpAdDSPZVwcDKc64
kUp5SYFRooCD5of6ak086rLyQy5MkA1VXSDV3JCy1IwYV6NI8LdIynlXW2iEXktR
Az99kFrHCra1HB78aj7E9kEJFbIlQ8H8NKMtFMCOzlXkiwi21jTmwWOI3j0AdhVA
i0dUjEPI7hbzvnfdaqoOnpBQ0z4kIYne3zP1JnmZVT6LRsrc9Jpoa8rc2ihre3kG
619QYj74TWnrOU+/AzrnOEWw32acZjWPevP49C4huSae3UDkedhCjnYwDp75gcE/
aLWGYsE8kQmiZSRsCwC3SxT7XDRvdIMCu7slXU9Kbs8Iz9C8pEmJQRM2jFczkOdK
4kscaso0gPQGUZEMScHjygyxAkOkLcM3iqTy3RxNAqNCAZnzLBDIf6k8GO8PmZOr
6UpGh2zdboPwqbUGYD1HvBMNRPx8FGkEMhdja0rpG9AeENxr8lZ6l2BxYErAC1mh
LjEvEmEL3vMxWJ8NZjwZG1jpt/mMD1Md6zDMdR+FDL9vnvQd37kqHYPq2lb0+yeK
omtFXZ160JDgWwOX0vhulHspB2C/PmcBgJUIFM2gBjFiF3jrmb62tCdeYdDZ0Biz
UHm3TNYM4Wf73dYlvZDWtrsUqc88JMlvF6h1HT9NNlc0JRW/Bitu0lizPUV8yjRX
hkJ1Tyf4Ykcryo1YApJ4x+8ZL2lSDGfB5GtpraALxcZvL4D6mmA9/2TtYP6y8nHu
rB2xDYjF8iG2mPobqQuJOsLRhRXLyV4faDvLOWvJLKTE5hQwjZ+hWfenjlal3vph
95PKTSZiqnwXBdv66gDlwaFBswKANgeYHSQbsR8JugCUBZDFe6Zk53R4Hkw+PQaN
+/n8cRRpIUm8GcGJFZZK+hwNaqJAjI6mg337iG0ud5WMztEEV/kT6WmqE1PRvbrg
ZGiC63ins87v/VceEOEiB+y0JZIlUtkRxideGy3lfhQEQFC3e4Wib0/I/PiOfi/1
cOi9jdT6LfDTiokF/ArDcRHXnJoDP8Rn3jJljwBqgqenC9ECRpwbrsIA+w3PZar3
RSf3dnc8Dwoth26OcQ979EqGOh5krhLb08r37i2YKRzjvatZiyQHvv+CE4Tt8BjM
6YHrIf8pSr9GKibGJ7ev0+sCyUEZ7UvO/7zEPWiqie0W7k9kkE7UQuBq/wnh3cnZ
IepKqnKOSM7299QZJsB+ReRhwjwriTpsiRbs6N68XJPj4TxPdfQDipETUWPy6zi8
X3vI21P/GCHavvno8qwLoyUGQLG81AeKqTN3GakCqgMlVZfXVcsqCf5XBUHs1tVJ
GoM3Q2l1QbfmrXKVsEwxUg7apSp/Sb/Z5VkMghf6ZXA4l0o+uf3COLZMsJytjh2x
j6o90FLfNmgnrFkFN/CnR7D1DEtdrnQcIhIGK049zmPgIc5XL7BRsTA/676br0fZ
FIzQN9txifve0//WWV0KC4nd+vfFswDXMn/g2O9y4Wm6SB5LbTq+KPlloqcEAQhd
3gARSbT1VtN5WZa+KkK7REsXN3t7jOSB8lnsulswrU3gjocPDu0/KiF7N9tXoB6o
CCU1KUILlCjn9XKiQd+PE9MDty1RM2PttAIDDipLT0mTYtdOuyqcZW71q7fn6baY
hV0ZsoqOrJzMrPUInoM4F1SCTiCKQmpMeXTOpJYV9ueXQbFN7yPJeR+7mylBRkVO
azOdsC47L59vlkCwvfBTDeFKYeKcKanZd1kd4OmmWhWgyFsvTtVUhRcArMag2LwN
tYwcdXrNJlrlHI4Urq/fxwJ71IeMKIdnflzhm9jVtc0DfF7FYFOFHdUI1MOkz4Ke
0Ocqf/9ItBmm0P5oOofopBO7JnYooGZzOnK4T3YqkxFS6LE9z2KMkBrk+5TfleL1
/bwo0m+viCRd1b1O1YMvGYm7iCu0nff3R4TRdJ3zhdHeGhflfAUIo7Ntr35dWNEW
q1W29o5sR2zhuwR+hb+B5O2ohundiMVy2M8xsVruhDodKiNupSBt4D2PDjhGOvka
JExuFULIvp3baz+nQcn9Hl7Fn7g+A6cZ1Nu8RxMyTq6ohVHWejAfg0RAu4I23dwo
dJ3XQ5qb/hGfyn6hzSq0WFrhNkSYyc7GBZ0ozJLH399OlxyEfxMe2VMACjf8JI03
cHNtRa6ZpMDLtLXuKsbJpVIbfvJ76r9JnYtkFpzmepHRX2dWuLpmT8GkegS/nc5f
BBbg/2KxyMpSJ1PjOUgkctq0FTlUTAAPNERH+yBnchL4EbjZP8cxkbDWjww5thhL
SvLJsZgdu/Y4nmCu9WrZR/BiAizLqPVFAiL/I6RyIX2a8Yt8+CmRRHfnRxa9KOtu
mnq/FbODXHLZ9C5D5qoET6ZNRJCFG5yyJNr9N36pxQ5+SH5b5S5U873FouSM50VA
V4kG1BtmAf2EVqYJ5Zdy8A4Or+wYc8ab7eU9u5nKH5FTuDGins4+/ot4BLWJB3Ay
lJT7hf8l5ZJE2NVuOCb3af1U4sKU0CltYoSjdXSCOdC1SbczTXKjFqRPQOOR3Hvj
xBk+nRVrtymlc13SLCbLKt2MbCtcSwcVX0G7VFX3TcTf03BcEjdA4PJvBwdEy2kj
8EFTstXvVL+nfCpJ6iH2nLxPSyconCuNTsfSxNYKfz/3PzwkqkrQIIucTLTdncwz
BCfjdHU+hhjLpZXisKaNadu8ef9GkkmJDUyGAGEVrW5LlQlX9heAn1kjqNK4pqNB
6Yiq2GN41irngwCQ1C08Wk3yAQOCGrQwWVR5p9Y/Waw54Fu4h6bGg+rFbgrRYnt9
GNz63vBxwUs2MmOg2emwnOZ2VZ10q7HEaYExOfjMDHn/KnU127uuKSeL5OINISEb
EsH1C+ZYLdSCrjR9fNHu/E4Fko/kJcCH6F2vIKMfP5ziwoDrOrV1XbXVg9sGsPKb
RQCoEbkyVxFl99DjsXSa5b+aMgAYevAxuu4uw6DriWkMc19qnrtbJHX8lWsHA1Xd
gjxCkQt+dkJAxXGnnsYQSEonMp9IoHJOM9hz8Kr4lrvozNN6sx4p/lwJJJm2nWA+
veiKqWxwmtTSmYo9FcKMn1vNRI9jpK64MGvWAC/Q7vN55mfewbcYUkn26WVJM7sd
ZAV0I53daicEycMGy4BoyRySB84hjKCzWRFbw5fToBDmbFBcREEVp3X3YPrPa+dq
/ywg956hiIT+Xsk0AmELTl6NjbrsdOfdVxiD0JFw/wiD4J89XoGqQabXI/qUBKx2
mAMwSP+ZU2iQXCz5/yQnx/gXEUqihBPKmH3JvEuLc4uaAADCufYAuR5s0vNtU+bT
mH2J6UER5ng7EPSC+/3FJU1eqzh3yKHE03fUhgYVghZE1LgKsIJVafh0NubOmh8O
gL1znk6rAALPKrEsd6Ns2ervcg6LF3vECCAqqTIsUygeyTD7zocS/mSXIsrJTHE3
FqxFm/so0SZyOUTeeTk0b5j8JSwB7/xjgyYpAuWt4EaU0D4usTxorC+u76ZuT5zw
0yJBTqROxfbE9ewR11q3tnlJ3DuohnClD1Mc47BimtUHi356UMao3oA4+L32+TuB
PLkGfjUEr59X+zNq17z1RdnZhg4fFBH6/a790sSXPnn3Bp7qzOG4lBdeErfWovQ9
wzmTiuyUBcPdA3IsbWdw+qu0SB4hxNo0e5dWhgrNxVpM9LWh09k1yqhkw8g3Jdhc
bfR4FbFVTTo/KUgm8N4AjLrs0q8P4Ma2UDTzUpvkHbxrzhCbkGHeuJII0bW1zgQu
M4Y0dOb3O+a84J9ejU7Yehj2/M5qqpU1fHjHw54dJsWFuPgB274jq0sJIaiQXxUO
FeDEhPQ8Hs/CqTSEJzktbTAsgwITPGfX53soBo2ogqGkwMdphpc1SF5ziPTLbcUk
wUUyyNjb2Oi5aUFfFJf4qciZ0t7mf+fqFWysWKG1Bpma+LzvQ/XZ5zCR1roNCmXR
HH70P/muUhkrUEErjGHEHR70tYsIq5G6zr6gnDhkWOfwTOQJ7b8cn1lmir0IY7LG
XhXDoXnrPGVnvMMGEV7wWaHiixNqoz4ZUV9g3JOIU8nYYtAw9G+qBVV2NCuARjTB
xu5+mleINUOVaCgXWrMvdXhR0ehll4k47svQd9xH2csnkQNEMKbS+nEfChXArHd4
3gm9BcOyJGe8n+TrfCZsHE2RpT6m/TWigFoVTxiIA9AZdzIAeEPz41g9vGICi4Dq
pe8P9ucIYcznWDA7U+GtGg55ne4Xbv0CyE/njQVguxXc/llRiy5r9mtVB2HUwQlL
pYrXoyBgAwIDMUUuSdpqVgqF+hUhY18UoacT2e2mglw7iXMfszATnIIhlK1WaYDJ
2b3IP1L58qxGRNntFPD4ERQ/B7pEtFlO+cefOH4x1SMZiHaxYww7aYQasOWl/Y4z
2VXK3BR9n8IZSOXT+A8MAI5eHff5DgP1CaxB8nfYwM2krrsC0rgvwKnDg4+3ihiZ
qwhs3sf6uc9pk2vpJX8sLNmG/K9QzHFb3y1tU9VePWjt5mbuSmT0oAo5xMGonPZp
dvNJ/zAYKCkGY+QVUgN+QecjqmB8mgzMv3JRANGK1j7qdyKta7AAQtTk4QckBnQN
C+rAg2b/De6g3YxL0ECJjXV7Eh5wfabRWlhmndiV7wDWusb3H0mA+SN+E9AoBMJG
rnYHybW3+EEakv7dyRR2GFcb4iEta+2+rSCyvuSyrRtDu8Df4hwizUDgicDBVJV2
pmEGaJWU5psM+itZVsxYgJ0Pj+YmzLmArjHOKZa9gHM6sFK/obc9n8rVJfV2vbwB
utLgIdPugOVLNFdCHYUD6la2oeK8N+QY3VbCFBJNX7ci8xGn0A+01IkUE6WohX+4
sKAzOm5sPCsf9gIt2XXdBVIL104ICy2wRmVUIhqtOMw1nWq8iBYflBJL+YDRCSMc
rstFv84ZkVWYi22K2Rdt+1qq+aD5NzoIbKj7mkcGZ+cSSDrvcpuEZty2tPbMAzzW
N1jZoW2UQkooTEusn1OA6Cw/mmPZ9pLBB99xd9L5Q6pmhNnn/mnjWGDO1N20qOio
zMuC6cUriPqFiFA2VjlhwhC9m6vghtcnXjVKnWsjI9gDAgQJ2mPDD7qvBpSf5OWh
1fG8zlA/dpJJz6kv/etmvnrxIelwqhsP2muHlBOJzTe109BA9C/bn3mores5U8ZY
TItfx1VPFzW37kz28dTGKvHCvkIWDTsO0dWwLLqnoGDy5Ftt8Q8kqp7FDx08BcZt
tXvlknosEOGBbdOEOMXYhi2hLSC1vvv8+JeyHEeHaHpK0qpCTo7sQQWI62ZCIwZN
Y/pz/HXo+gI3oqhQcNn8yMBSjcdz5H6zA5N8zs6L7fX28qcl9mdXk3qgN3YvDPct
Da6+w2pnYZeuVwyLiRmfEaWAtErPCt0jJO36OsuU076KtboH2yQETfT6kt3cRON0
y+YJa1WjKZYtz+g6lX77ZUhUkbAGO95lAddDaBGDmcrrSJX/gk1gB8LwFvC1GRFX
uU2H93mNTSB41rxcfOXeoI7QlbnSvRFLZ/QrEu/r0ZJNcsZgUeOFUUF8AeIBLqGn
dR2mIir+ZhFCKBB98RqXP5uL7khN/fAnZAYJ6ljJfEEfS+CaSW93l+l8RJ6AR7F7
0sGXtVTSkTw5Kh3/lpsFrGjwLg6HqRXIyQGTyCEbCpr4K8RN+EbmFI+IOOgtAH4w
7kQGj94l8bVS0NlzbK/YCVieyAhJ0dSw9TxJx+8xQvTYN6KzknAhG0TF3QEW8oBz
F+ucPO6OSY9d3bOOLeKHHwXpCLSpg6QmPIiL2lQA+LdM12mavEvkwBnHo0uwiO0S
nNrA2AHDse4jbvA/trHl0vyvtBOTYk9myOOTX9oWRCLYZqWdohwE1Zzt1RMaeHCd
S6Muff7d9+Rc8Ple6x0h4PGKB4hGHRs3sP6KKsLowrsyD2Bmu3yN5W1onwuxT7Ic
mz7OSjdD8RFq2QXaQcKb8qE+4/ntNiecKYWdaLaVSlyMbm+Carq8M9ACTkPxyUMQ
vIo7uGiC4+4s7uezf4dPUzgJvY1zlcldiTn5Fu6mbRfbhLRcbv08BitRmui0C4Kw
WBhF9tBTs4i8XPNk5urroqSIX3fp0nJ7B6e7jl/TsBRsJJrJW1C00AbdlsJ9jy7I
ltOlh4N1P8X/TWKeL+e79FNoGcjDX7SaRPsQhAGL+pX6IKYWhhlqruPafE/z9yfW
p0hHKNf8L1fDg6/EN9HsUZMAQbxO33Pgb9FqKaZw43Eo+0UpKUHBcUsehfjiBpRY
OZqrvl2dumphrNdnHKPNt6cmymduExmJ/KZxJiKkXaHQ2cuCstX5d1B9qukWlXg0
vLSjgV1NKvDMtuoaEeuNCWGEWYmgCuMEMM9CN3lI9bYJ5X2lNu/UI04xC3WNL42q
ZmsFn846f9Tnl0d0X2tIL7Gv7CPI2NHBtNv8+GEVpKXfYaRh7nz0htVJntfkCwX9
JRrzS3WbDlrRgRTbUZBJy2cT3Uzam2YLLnS9ibohsd1LIlbVTPfJsDWpjYXaWJ4H
vEuHpheXUv+wE01mi9Keft6UJ9v3AlcBM8E3XqfkM5/00ItR5Kcn7wGmW8CFvZFF
aC5YjhVuiEjNEK1nEcuar4wWKGpg042Q4fPbusKZjQiRlcH7Sx5yiFJxorZoJTCE
ZJNSRk5stjsvO8ZlyvLZq9APmMgB11Dyubzo6fXWlctMOydIdUMz8AZ/owq7YTng
E4sqXdUNp4Zb2k2ORE5C9jpHzIFSAcL96EqfLLzbLVWEiOCGvxW6hzeQ8kMRfuDq
tM2PATbhM9FhLSnEOY3vVe5c0Jpam+e2o0WApMMOauMYTm96uAe0wIwxMqKtlwNn
3tPFdSIx329mWzBKPhVCbugzkaNWzkzLXUwUHeMx8ySgDpkslNTQe4OjEMixRVdA
f3AXV3MGr7r1J/6wRZ13z+FtdTeIzyO12e29YN8hs4Xn5Cz74c4Pj7U4ZoEXtLjI
NvaLE6tSNlbc+PuIrD8bOliQX/nl6hJHAQ7hJ6XIQWJ+M32lq1JHyVdmor4M5cgD
3g5ZwhJvlQsHwhSk4NgKZdLm2VOYqUtybJzObPcBYlm/uV9eSkoraC2nVj6dGeJr
5NcReigox5cGAooZKei1MqLyNXuZTgOypC/CLx3GDw71I7j3MiFOXkfSFxh+bVZf
MbtMHRMcHNV+rg6rKod0042pMWv39FH9IHeiKZEHxQ8=
`protect END_PROTECTED
