`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MeL7QM6hj53bdoeJ3Zm7OrRQAaBFdCebeN/9VL9Hv6eZWdEv1B2hwkS7Rv/ORQCK
UdmnyMnaUhwe7q0h/YEgue65HlzaHKhky33z6pq0GdWdtQXdsT3XpNS+DAAxYE+u
6YF72zHEcVUtI6iVNdQbmMTPjCmGd77SE1k3qfgPEJqkx4fJTiz9dftBt7Jgp20c
MZjXwxAwo/a20OLIZIZTh/V5Pv9MD76y7qsZCoY5hcQNUdmGC870lo9KKyGlXI8P
OKuTeQxzgTzYlQoUOhaRwd78xjal0RfxJTuaAQ2s7Zvv3e5zg0Khaq3MYxTsLRNS
goUYHoE2XJ2RGSt3XBTI0yyBnI/POwUFMwITvhLHOzU+BW5yMacg697cmi9806+g
Tko7H5tL/qUomYlPnDe+3k5xE8U2hPBWz9bv6jb1GF0AKg5XoC2s8lB+WGigdAxo
bfv++Efb0cGP7e0cI8j3EN4mvEJBHLvToL1I2gMbr80cFyeuFku5DayS57jDWezo
1PfklH1+spFVkBpcqhVu40nXGkV3w1ZhW1+eJ5fk4KcDTp4BN9lFvs0za0X8n5CM
b4mBbBzLKY2EGIx2fAj7SfiBckvasl+2TuU2jD06ylLsiqEdLPozHCSA5YRTz5q9
xFRpjvX5YscWR6KaD3/qFRzCRrIfi7xrmBXWaMbWdMTUTyWPMO/V58R5dVrGo4ZD
PkXlFDe6kfolZzeOdtj05GcUupjpOITyApTNmVIh2MtW4hukHZXNwQ9l/4BakdKB
iFCEnYwoPs3GwmRGkAGrWizmxO47na5j+dOIFWJA3kdESbZ9vorDBh7r8EDjxkfj
5Pd5Csu1sl3zZQierpTd8Gms/UfHC31gs5JJLlhwvPzejDreyDfEsF5pNj7r68Lk
E+bCE1gbMQpC/CaneCMdPK9JR3+aJT6Hlxj3hM8xUr+cMDQA5cti1vOJitzKEYSJ
72IhXOLqyJWV+cXgThWzp9rgXknXNESDZDXrq9GqRUCeQPUJ0qFUeJ76b1I4oM7S
PmJladpo7h04q5A/cQQapRvux5r1P0RjsHWtNKy8puElgta3sz1OCLIy+N8CsCRh
tva7F2wX+f3dhrVAruNdKRFMeW4CbmJHqGwOBBS61GhYLaxVlyRH7iRAD7Tg+r/n
YF4AlhBtYD7hAxMScVwYeCq6ibquKxGDL5r0RSE28HL4fULmD5dq5Z2w5y4c5Rbb
0i0pjgIc7+7uLZa0W/ZHW5u8y0zqNWpWK5Oxw9RKy29ltlXRhRDN9ViN2YMx3cOo
a/Tpf6Bdu4ZYi+xqUmF59njuvrNC3lSDE00wK0H7OKBWTvy+ZaykSU0YpwQfoLDc
o4zWlXZEpGgZ2pXAKdML2eukHZnJoaAGvOnwXqw057/CIuKoTndishtqgY8qGjpM
MyTasPb50YfqBFd6FjavmIk/rY5zwfPNdVU8UjABmY2S9zItvZs1/asm14LCLNge
7QtM30QmHAFDakii5iJPJxoO954NP9Z8mr0qxV8hbKblGsAzDfwwf2hOMy4hx6Rc
LuobulrNlTtnoJVGfSdTAL2mcTGMT0QN8e8Vplne2PkY4If4BRxhOF9P/KUCry0b
y1xPjnPeclK5fxWtUh4JeUsS9hZc0mExl2EWmpcYqS1FkhADvdq8f1MBFhvPBctw
RfoJJtKnnWwkE1gH4Y6HYR+lAC8BoSVw8woHlNqodAoyJHID+25/C2QL62uhrmfm
k79oiQ3MWeNbSwemRWkQJwaLea/tp6flz48jQQ8dOTw2+nFHasaWEDfkJr4JuB2N
vuAXjYXI6cxE/U1lU10mTzY5fkR/Z+2PpQ3oQiWpM83WrcxlpcLyKaSy37sRd5mo
1VfOVap/jnY7jlkLLUqhlGjfTtlov+bYQCvQ2/TspzbTGJq7gdgxQT67dHlJBg4S
b7npqwyap1T4atLe5d/q0E+wlJbPxZX8mgOTga7e1eFUlaoK6Q9elWQi+hRIJn2T
3G61C/7XZBYAa29u0vRZuDM+Uy8MFPt7m8BvmxveTx5uXDmNQl01Cc7UiCr5PfFI
HVh4kExIkh8cICWiUpof59CLiZltDK+J+pkih+b7628bPyTufsBLzM0hL3milMIA
/j+tBot8w0xmW62u17pGi/lU7sBDl5j5ShEek5G8OV4KWYX5rKyAIPI4azwTHVWN
QuFtG4LL7U+71GOVxvj+eGN1DPGTcf0UqE4ps40hur/O5t869QbxVTItrZYK4bKm
1CFV+Fwpp3cU4jAQjnPp/R0LPC1nH7EhvlrOFU5vZV2ngUBuYCQVWgMkqdqx9Q5l
q47GAH8+woFFVgQ1XIUYilgKDesmSCLRnHGxLqA9f0EbSPrvtQGN2H4FVgJ7KbTq
3sjHAgl+uxvA/w3chdtjXd4WOYwlQFERh/7CUBp+2G32tXfUOtqESPWY23+ELeLl
QdfyJMRyr4DNZBYbWUTwWt3KxRkaVLm4cltsnMRk1DW2MVtWGTumkX2fM3KXVcTA
U9VMQqrRIUn/5dYedthvN7V5sZsoS1voMxd10/Oy6ikWwvViB6JOfu1LFPATyvxU
kQrhkiaaj2TAhfqj7z2C6iU2rrAsTdmnPOlIpoeQD1o5L/yayv/T7NJAPCJG8KlH
7hSpnFFVSuUnxaogm3196hyv/2fYRcYmAzeIV50zt+xoM8VU5gOGdpRO9Q1UZ6Ub
p83JUaQY86AfDSf/CTmMt0T85jH9K+0rFgob2MCzGpebcBqtffs23mqIrioIEvjY
iMwIl9/lrQruKNphN4woNtbK6UzqOvM2vsYV7gcz3whk20h981A7ahUIQd+i6u67
k1gZ5SQwzsA7W+6e7BkRE3hkz2AveqdIf3FyG6cJNgxBSAJsjXjy1SDEOGjEC1aD
0pZUkE45RreN96gxnVqbMoj5nKHlzvzbaaEDV8qZPdVOPdTHB4kmZC09gfiMHJXX
+TrZaqg6q0l+aQsKWcbaKOMAN7xvMebR8Zt6kzzupHgdCiofans82ICmWe1iYk26
MwKoVZ1owRAMbZ2XxBqa8eKGB4yPv62KAYKN5XmBD7Ge8k3d91nv5WWhwsf51pKV
cJQAtFK3Cywa0RQfu/g5VBS0ato/FMeKAparL5bhnv+94/rDIMavSxp0meHhdV7+
yZC2lOUgXpDr9N5ZUWb6SQfJiwsEpo7C9dp55KBE/EHPhGAr/NX0+7ycCHV9GyI7
Bh+pXULSP/bsX8o5JIIkH7MAo6ZF8rlyGcPkG4bhLwrCT/CHGoQ5Pa2YekHkfgvi
RGS/cBV9oVVQ1uw4u1FpJE9gXtEt28r8Py+E3rMtyfi6/1f3oVPt9d/V0Gu8tIUs
kjOlNN6ADXWQWpVj+V9006+uJnfu14ZtQZFcNh/+SEyuF7bsAehdoQeUSIwc1hGX
PByvLOZvAhOMQyIvyx5exiaelV1YpGs3zNeTdtdYEsnzIYtCjbAXt2gGIl+gNSd+
VSeAXxIyzLjMgvifUVyQUMJOsMwxPy0NC0ghZilb1V2iMuEK1T3VYazwwuBID6gm
QXKf18+XwVL29mzLZCLwfV2RpU/cjQISjg/YQdfvJPDvww2h2msU2xTR4TKgo9jy
RHK3LVI+f2plgWDTDAJq8XMOaXY6WoVDNnWhUh6XVaVXYaIz4grOmFUEC/Nx2zIh
9bXOsZ5xySG1fclbMIW3/UpyqjDmljLkAMJMeyfhp8k/Dmvie84mBL+lI4O0lQPB
N0NwTetEHShuM0BC+fGqkdaJ9HpMKBwCGPjtBLnkU7j4KVTv3ZO9gUXgipRMbqYN
gKc5LNwKwDI6Jjd9F+iw4b+z9SW4bECLeEeL+yC/M433LoY5vr6qjbMqjU3wwbKp
IUGNWWRSraoej0zleCH/MzFRu/pSVfo4GAsA1LjAoPAjIp4NMaxOEeuUZZOtoeH2
JTULc7mLiECR+OXz9kxJPDIgG2KblHDMnejKfYgKqY1/Un5D/AX89nekMIsL6iq+
K3KjuRLim8dvOeLIV43bnWq3vw/o5UPXV6GokXbIGOnsOjfJawlS+i489zyjXToX
R6wmm/restgH9L0XQPZJnsH9uSFHVuknkgVuWknYMydlaJTAHGd9dE+5L6KLy1N7
e8MlswlFrV/EccpukjmbwJs4k3Cexi+UmNI9S3R9hvM/kdOBeAdyHnXwNUUUaXcr
kg4wWEym/k4vOYQaKsqzZHhWGRyc3ZJVqdACIG2sUeGIiSeHaDe3DgcyO5rqo8QE
aKAFYYwtIzYpm5+0mEwQ5Kk83PsrEwZhfcY61s9XXWlIN7x09RdwNZAjFPYvce0X
ijrXoKDXepax1DtaK0ldVJ6hZ1KPJjPg1Mu4mpbEh0THHu9ATiiXoMcu2IGEnAIV
9s1ZJwZ0MuaKNfQLrT4I7d2iRhVJjZdqtzodcVAyJN5SxF5atEKXtRObhPz+QHq+
fbSDVL8XVM04E651NPuzPYD1/Bk+EmQTz/x99s7WPna0rKLG/h3Prpuj/w5Vvxn2
PAEluezIabJrgE4XLHNGlb45T7KbRcc/O8j4ns26O8Qqg33NHMwjBDCFxpS7uOZa
lX+NLyVmgQkD5kuCdEmMiLxFZTEqf1K1q8yxYgtdrrZzV8ltd2WmflMa1F0tHovP
6/Twahp5Lb6VmcVrWH/eTrex4fhLSoSAx8rN0+Qtsm1HFTGglKf3x2dn3a/NilCd
RBhdQx6pIigCeUW+KQYqFLv7QQUZZCYfPhmUOIa5Ke52wx4YynbLnJ3I3KfBF7iv
R9U180zI8m5fcnaM80eXBrqhFgTB3llRy+2nAEtaSAT38Z4/XUFC2TQ8/dfcRNPl
hUQn0HRA+oCSVciu8rpz3nKtnC1spfcVsv2FxaTTz3VdXyGGnTIfuu8fnUwrMw3j
0tke+c2vuAygvfiregsFJeh88feZ5pHPdJ/mroXHmhSPmjFFTmLAq8GlBPhKja3w
p1iFyU2y6D4A/7t55dCiOZY8hmTKkdlr4oP70YOJXh15qlkZeC37ontYboL1eFzh
uqA4bcvN/ge7/uMBnV62U74HPkOaT3KlM4WjE75Z7Oa13qVsUl/SvPqmNqijHLt+
aDE76yRbccQH3ptdUyzAGgUIROGDVtem5JBoBohZO/Xe6cR8vLvGn9/GLUMmml+H
4XEcEnWckLVYW++0PNA1TJ02crTWffcdpGw5nTTz6qCz7pwgE9XucEqKjTmuAnQg
9mN6BJbWqleJ9LjrxDz8GqMfrai+RCw/Be5SqjtsM8zmHqYV0vq5fmHGmAcP6gPl
vbwsJKICb4xx+bxGX2ED/pd1B5EE53jKK5QB9fosEoiDqx8d4iCfhBD5687t6GCj
9W3dxqZ/oK5BPC3+Jr4gN9Gisk+LYmlc8f9cFbwFP8bT57uZaQ3QxFGgCg5Xu2dO
qbwmEKl+wECGrrR969m6Ioq4/ZomxCf87SZH2Y0LjMqKz2KiYn0P8V80WjSCe9Dx
q/hpD7yOGP/N3BZ0+94zSxAiEBGfYDsXJ14BnSjq5/gSHZCZmwZI5Um2E4A06EPR
O5eXIZmVzj3Ib9RnPWvraVO/o+Zm3n9OzjICkjURmTiOGV8mDvFIewvOkItNhGca
Z79v9ukPhtvUmiNN1VqHLaWERwXAgmut58Bzto2OxD9MjdfbQBTVlXOsQ1gfglxb
wyRq+5CQk6EYRiOmQwd8Hc7P4sgzcCH9w2mw6409i9/VKdPWowtaKQvf9F56nMvr
G94XfDFZ9XbAfLF8BooHTPTAAzrrzVqYk/PEbJ/j+k+Cww/8t4GkHb22GfHzgWgV
KLJmav8VYJKXX+aI0cZk5/TjufB42kS6/jb5T/uRnnIRA1RWhp+DuBB2DvUaD7h7
vWtltGXh5SrIwrYY6wcSXmW0dpw59HTGsWgx56AQJDFv/en/rwz+uUSkrmzm5g+6
dON4kbUKo1mB9T3u0H0sgtIF5gtQy9WGmRtJzdCuNIpLi9di9JFQ5zRukKeJSStW
JKld+TacyzCA0EFKjhd5tfWJRSFUz6aHF34yxfFq9noLJNoulwt6CGvZTS/V18YY
41m602y6a9R5p63eGTxXHHc2U/rQ378/HAwey3yr2/wxu2YbX3ZSWvNNtgfG+vNr
QlXExcUxJVbv1/zB6rEdPze27hMrM/148tKcQVetXz8XAmU1ZYO8HPC+gyrrWvld
TOYWF6aDvZdg+PBL3N3Mp7hIsiie11jT75TA9fIVcaJjMfbAH65pmxCXO1CHx+Vm
Cvyr+gFLTWi3+R/ChBSXHFNmse9MdI1MgOgr6lu3Y0jyOqkqtchE4wdYMaKNSMoU
2yix92TYPw1/HZCu1yNpnm3yoh1JlzYKjBPJE1xwVAEZxx43BTD0KSdv2f2od4HS
5O2ELZV5De6iFSoP7mZpzXAh2cjU8loQsQfabjE6c1exG2eQaX68LiWcis+GGCHY
GyFZGFUEvkqJ8bVBMZyusO3p9tKU6S7wEHD9cchytc34UszcOszPzsPifMEa1KcY
Qop46FrbmypNK0RQtlDVAAmVHOcbM19Brpk/Zlc1/aEvibSlXe90TAs3YSD0dPx2
L5y0QPIHU4aWVmUUPvjaaWFA1UYCRDj4H6b3qa75JudDH3wi25Ku+TTrUGKFpKDd
pJlgtViZdSfTx4kM5RvBrkran1cpZE2hqUEShFzKyMCOdG0psphquotMYeu511lr
WGvOjmHiJMEQH3kQz9Qx4SobphMoLslCgu8rRPjqbVwIOwZbA1qsZSXKMzOy/qr4
51XgRKj3w/Of+0i+17nBcZlP+ZELi+oa5BHpBEA6HxMVqdQrk6TBqM/QbFIg57nU
tW4qBa52TY0tseTFmNxH/hTV+h/gft679qqzIb6AUgZ5eQ5NfjeFHKDEKRvHNOTH
uwNzB4k0QqNXidnds1/De8xTT8b/D74gCCbNvxMuWa+Z63tIyT6KRqlHo/cUhR7t
WvJS/TGBE7s/PnoeGwiFc8DTTDdXLG1WtoYEWZtkboc30eg74yqetS/rhLFBvhk4
oS3C1LJuIxjF6pj8GafB8uaYLTBlE+aX97fDvNTxoBnXt8o/GUSXvBS+z8TRXI41
iYBAMqk63+aDIuNQIg1MJvZLS0ai2MXom+/aBxtb3O7KHJ4ssI61W8n77suzK8JX
EYwkJYOdFy3mqjpPGepLMwqJDXxF62liH7aC8rwI6eAbXGgvJxjRFqGiv6LR0+or
WZ0Q36C/1Arum0TR2IGTAzBtc1XJ+Fjuic7xymaJqa3H44lX8JvARtVLYc4E7A7n
2rXQ9oydNFRq/bGik0bfp2lfsXpw6h41eCs6revWTGXQnTlI2mti1orJlMIW5Dzf
UieY0dgztA9x7PDzBMGznq+5DSYf46ixY+7XaPX9AV9JXAt1Ye6/WjjtZI7GShc1
mFlPryKDL9SLZwBaG4WtuNO1TUjTn39TEXGBGzwOk31okqDxJW3cPzvdAfFBoC/K
yKKzk1OM4ukDevrq5jG9Vi6jfqDcHHcI9ec7FajLHNAcxsRFq7QpLCSmlLx7rRU+
GcWas8kfl3+1pRojlym8cFzoDpHfsrcO+ed8pirD7pl87cA4wtDl9Q4LjsR9M/hQ
vDTHBrV575XJWlD3iIAS50j4qKpDm8gHXv0aeKtVcladfcCDquBH7VAeNWiyrfmY
A9xtLury688UHE9QtHXCybEtNPeOr1yA5nJ2quxDUKkXirWIr1cm6wwGrI6JzN1c
+yOuHd7xSnmI9visRQU8gJHniShV+8qGUVBeHcFZaEmxJZVqtZR5hQzItUeqxbG1
UoC6xDZHkkMME//pQ34CmNRy0KG5r+ms+SQKrw/hBMSmg34pSA0krdlb7zrTXTC7
xrUH3zJkEyHI2FcPFrhYFY+nFgTyZtt13iZV7zs2/qkywYiK1P0tN8bXLoN+FKIJ
jaBE96Ars1p20roq0ti3JI56HdpMj3cx6kk4BIn/oZ5yCZ5S1oMCO/FsX1fR5AFQ
NdJ1G4viD31G8LWV55HnCGFwe0zDIVdm+7I1NLpGD0AIO7Db4xDpzOKraMuZYqml
i9OR6dt8Zr8+bid5qvdL05fbmWeSsCeUAf5pY4pos4CIWpqwA94YExMK8IHar2+2
0hFI5GnLbWwVQI6U47zdciJq20eGVrP8MHZ7zYhUeZH+33lgh+vQsq6Zh6wsLzBm
9ibFCEBbJE3Sjb+fP/E6sD1e/aHpQbObOJUnB7DtGSDO4ITFnuL23psv6/nRzVZ+
wXSybFddicnxb+Rro7MHYuOoQn5bGXJJxk1/qhBfsYJQzHiP+d0/KPTAc4B7pMvU
EmnXrqrzyPzvLBDwVIhAX4b3yVN9xZuixm/l7jcO/P27G5/aj4DzFl4ze08tkkf8
/U+bJtevPARVCP9oSDtYMkegWJYNEfqtTUwjn8jFWwnkN6fSw2tUQzbocS3ANKAl
MT85Q/INqM+6ulXKhMPMl4l+g1YF/rLGkRyTrWfWsu9HJqaQ5dG8MBoS5Ir83AdM
YDBv0Bwp1Tr3AzCNLaClIulnsLD4PGS8GpJpc915O/0iKYI14YuPSrc06gUka04a
Lb4KEHzWGxk2D5/zus8SHGOrk35k81ZJSYJC7OLH/jnwXCRzwRHVPau6SSl8FHKk
wVp4rWxhfSWc+2RMxTUC0wCH8br2e+u4TRLVfeSwxdLHNGXGu8bdWZvkWv07Uulo
mizLkBDPPFwjNvujbmtvvbxK7jUECEVglgNkDjePXO7v7tObJXAuBJRvrS/u2W3Z
OEx0jnlmC/pwUir+xpMsaZwpCNyaIeEFQqiwS8A4zcd/owuiBUtLGJtcL/arkDtl
kRBXW3wXCCIQLMu/205geZs2eexAa2tdV5DZsYHrhCML7X0mc7A82fIGy06GkUCP
VBOARXPPiCfDuRB8hbFdYwrH9T0jmGfhG0sIeRQHfrKauYdq6BVz6ZBpHn4ssXxq
MaywAdCNFWSBzeLpZhN52G6X35p5aDc1URCMqj4xJ9kZuw1lvpXMuP4KjSEl2O4o
J7CqY6jc7Ln+rQxjM90G3N3KFWteMMNOeydjEvwCadssIOUdsjPnftccChQqO+Te
acW6ukurO1scQaHQXhoFImYlhZn/VYvVYAGmHD7XZrL5dOBCVvayi9lg6oYZDq6C
89Ljw1UOETxE3XcLWsLdHbch9mFoRv5EBf+2zHwCiFfNj6HcWIf9t3tm8Q9aTioY
4uoEdG41rDnpJwuOrKB2oDJs8CPq/k+jGYM2sxBMSw9BAH/ICsZBhl4chA3vhdh5
aQvsjfDmulhrcKgJyXStQdSNrzPFjONHP4BEDi97CQc17/GEml3039iMXfocyu1I
A6Bl8LMHH9zP78o5nTAnablt6VxRzNCqnGE/nOKte1mByWHupOCilW/aLIO5UqNg
rMabi7dgGd7pNAxE+EG1zzp+Xr5dNLWUqxHGyQW+emv+aV77yNYn18LlKxDnqMoM
0Xcp6BPBXh74Dy3ObYzK1irP7tVl1ggIq7nP/7YGvIrycPWGLIOFgaHLrUv/SVqd
u+KdcU6aPOfTgz6o6e9GGPI/s5uGZVXrvyFatjOkQTeB65BcWltmZzw7WptfN/wp
01I4ewBWVGcMvu85JclFr9lJ9fIVUDpaAttxvT/rv8BVm5zHToJ5pxIr7uk9nXp5
Z+Jpnv73ERwMwKDKALiFsZI7C6uBUHZuFmFskff/rpGCo63ZUeJk17p0khgGolRY
ICvDIda+XblsejXM1eqUAQPP0ICiGqDpAL2isLxNyw0rjkXFCUSGP8TWfM5dc3tK
YCXD9+ioSYLR9/ymWUH9ccrtqh6xD9FvUoIDfKOC5aqsUuNeNzJiY1AN9J4nIA5k
gPOHwsufsAmST2LgUt6OLVTehKSsbC4CiLfYIMxdrxJEr3l9Hu4VIxWmsPH5yVdG
QloctLicRjh2pz79KFATmvIstFsxZXoFwQ4IBoNEOaziS5kmjaXNIpOiJ7Sw8Ydx
Ru3R3uN8X36P6sWFqLUqVl6ljzECtbs914CKjbh+QW+NzbD7jDBUH3WK8g2GvLoo
tuG9nBSanJEEkaNk+FbTvqOpJtDLZbcMcb8UOrvSpsIQURp6hZu1STT6JGiJScoi
irv7BxdIiegtMlQcgQt0qg3zh+B+7H1ksJnqbZgqE/9QHhzPLvONDBh2d77PVhU4
QSH1uZt4o40TSVn63QS4mVkO2Sk7Nmcy0I1BQoB/aovr8A6FmIVRzzeVRvCGlvyh
L5XFpUEkg4aFzlnY6ZufCbRmeHrNMg5CAtO00T4pWp0gcWVW5aCSJkvgj7DcY5v2
uS0oqjYf+ZGgpgHgeipt7klBmiHhHr8KXhX32VhEKMvUHkocXcLKB51d8EbcHQ+K
g+aMXIizPWFOhm21jLbL7hHFgQHiFLk5bgZcgsRZciAPna20/2hQrb1/YCmJThye
7zrYpxGZ+3HsD57Sb3MTzP7GBAABJN3EpvBvQjrUv3KcsIXhjt3R/IywTNamAN0Q
UHpQOJYgVnFDKy6Fsf9uLO7PjdjxqvcfoO7kjwyNT/E=
`protect END_PROTECTED
