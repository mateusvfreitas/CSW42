`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
E49TsWuEt7eKF9iZnV0OWE9rGlnUBjQWtLAlA5fh1NFyPN/l/8GxUcqrDYkXAiDz
BohVbZHI7xmQ7c577tC7v/RDmuB156ZSDpBzOCfmewpOK6VsjmEyYHAhq1ASBppz
6TfNQ2qjh91tzOeirE2iLAu9aVuHMuezdKgfdOiJhNFmigauYSmnqSRlXM2vxAV4
Q9R+67jBcvUPL3rbKAjasL8lv72eBMyp6xy7FzLZ5UZWY3o7t8HC3BqDMAlgKrWv
ECIRzNDTrNV8LjbyrwwwJFeq77I4poR5yfdjpKXJ4JVWkyeJZg3lzlsWKrD5GXzI
G2m1UUxcMdEoxbPEa+tv9e00PBekf3X+OuJ/EWx9dPB3LOqB6qUOS40xLSSagUOG
eU8Soz39JuAKS5k1coTdeL4IDKURo+SWph6739viuPd+G1bVsk0jvLHXYcXoCM0/
VVqSIWFev3acEUTKFy19zKm/+40aTmxX9VVOd2CLtLBoIjNL2TH0oOXC1tCARqQE
jIMKdcqIY7kcpoK+qZebkKoiOIMCfV6sFV+wKkXrNR/PtC5OxqzV3ZAqwqU2wivD
cVhmOPlGK332+X03OWaDGEZLuwSM6cqK271FEEA5ETMPDn8E8k2odYUgb3JHNpi3
gGLKDExBQJiAjEJ/5Pvq4YDgUKL+uaxmm1+wWG7ymBcIQBRx4EEpSLouRRLxs37N
jm+SIKi0YL8DBsErpCXhKsUMUuuhjq8WTdpv7geTDDXIpDTEJbVtWuBtxW07f5OT
llvvguYV4NyyHYObnbnwO59BBdj2do+trLuFJIhe+4IILlHvB8L6WpP/Ptd3z9W3
35dX/hcGwb3wOAOtEsqsmqHT/NL/dm4MsjKd5gMtUTqQXZg2vYXhNczNSTrHBT5R
x8vO+ZKD0jBKcGuUyteEinJGghVrju6S5GOMR5bU6Q8Cos8rktcC5ww7i4Cmb2kU
vtc2xaI6iNRQSJjoZfTKplFIh7gWaLNlqbDaRO4ltcqP7gM4wp7/9mhjt0WJEF73
Q7MpLfujj1XtMBieB1BD+0q0/hPlwp0dpY1GQrmF6a+XZ8IVrjsV2V7v9GzS4RLH
I6H6nan4pPpr0qerYZKCE96BY2piwocAve1+aI2fMYCdiH0L8rCreqkaPIxcXs10
nG1nSVR1ghhwWNomhhvp79cpx/3EGuYUigqD04tvZ515i+UagFaj+QUZtaUKc7tZ
VPwcWbWb6UmoDEu29trXhdes9jqtMLD34qrd9wMnV4cTj37lv0uFpLZLXQp1koa0
zjGI/IyLVSPivq0gDUzJfmE9LccrVRyW9VdTWLv2LWQ22iCnpbPB4BcA5yQXxIXe
kv3Or2qvKfR4KcuHIlPjsQSUhkabiWkNLFLf3gjekafSbdKIL1yz/smihaJ/4Hqs
aVhpDO7T56+bR+rrPQiC7y7FgjWmTjmIBurqqrpJyEMSFJEMjgeGMF5cX6T7BbwG
SKbbhJni6pIYZubV/DlNR3PGNM/nxtnEfqRTQpvBE/PrpeSIDf+cud8XDd/HnNNz
WPIRJ6G+siq8ggnheu8bJH1cS5iTE5jLrcRM46LATmyVj9m56I2Ns4d1Hpdhd46F
KhDs6lNE6X4LxwYfkc/6+Cbqem7QmjQYBJ26Cms7KEjrdQQxwzcJli1eVFThr2r/
fneRE5fC1rivWd8ekHZ8kSIFJEkgf12Kv1cwAITVvE1KckZSEIt++ZQ31xt2s775
MxPV2540ou269LRT7ZspoDlyyvQKqQsqOLQp0Uk4yfmcmIMHD+LipwcwpnAZAUfB
rnTYyVKpSOZizkd813yFx4HdKAHoFib0V8c/iSkVkWKe1TKuaUzD2Z4NcmWp7EKK
wDIsWXyKkhLn+VxFEgnA0znT2IVjJ/SvluI+4cKr76nvu8GkP8479n8dOzGPvwbc
zH6s+m7zse4rhkcifV0MZCKSism7rcijRqSwq1utza8n4pNDVP7DStuE1aNk2cLh
6RbHMO+LbL6vepauBhBuAg==
`protect END_PROTECTED
