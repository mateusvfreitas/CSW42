`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
/jzLsKh/nnh4miIU4hmncH1W0yjeEmFRa+7DODVX9Grm9XTiODIiD3Wm1caOj28Z
8mYCZS0zr7TI2gZTpmPCeVvC/lu8SybXeNt+toyCtChteSZE1ctRkoD+JHzWzcQf
jU02QcS0ZSDvttAfrYlu3+lsWwP6xWgp0Fx0JBCw3bq7PLKPnFLPH6fjyTs62v5I
cZ0J2mqDFJutqxUQ+HF0kUA7hb2ed7x/P0gVOuNNrdH33wUWHE7bDXVChQ+kzmPc
Zax59vWtJtHV17Oq9vhn9Rjnxa9Gq/JQph81putjCRPIOJGRAg1YDxrlgwNMBrca
5XRGn6/9H5MXYb/RvZBTLj0S6BlLDzzJyZPUOjdJZCQG7WnolKflsH2JtyTlI+UH
OcxrljFXU7ufyfIPFus+hnWg0Zu3HSJzlaZtBA1XUmmnivv14SSmwm2Ah90yyD5C
dP0vt3GWQeewHsym4IhW6/zaMyIJhWYsEmcs0YQozN8HURK1H5dorgkZTUxPnLUq
01Wbn58l+IfBkk0CW3CdLmMijNVC2y4GpKJYuo8+FcQzfMkNjbiqohliWBJ0zaOZ
eOSs+ApFWHzCZky68gAR8hoxhr8c/ceKueGZMjk0CvQJVdjc+enk84dV8e3tzLS2
y8GI3zZLPNlDbEBCJc1C4hOHur2SKUtH/GOyRfieJ4NfYYLXkI3UrOl3jJE9WRWX
n1FrSZGH2RDVx3gEQp7vYAoXVEk/spd69ZYTKPvsYpJiWRBilWuoAprZV48ITHSm
u9f+fcZSj7cWy1EefglPl2b8fLq39fBugyll/3jPKUyEdLdYjwkseLIpjlOJNTs7
3xNgM+aBFr4qGcETT4pUlkhSSFXpkLo8JdCNugttI9FnXZs6MYPOuLpPt8vU9YeD
RfK8vd/De+Fri36JJ/R7HwSN220a4eADstJGD4bw7r3SUCNxN1pY81QA4TLmxMUU
i2fug2UCEjAJqSZi/jK/t3gVbCXsoexiDOg/L3k7lQLBjDn5BIBiO9alFie6nDCc
ZY0Pt8bRngmbcPz6S9LhnbVTF/RId/vjw7725asjVhSaboEb+8aLJ6189vxnOG/+
gTnUB7ZVEt8zaUiVzbUdYEKiPyQt0c6U+aOUvz+X/6lI4eVS2eUmHm2YJwpHvwTO
MZfISrpHbLrax5NSSeU0sjoxTWgq5QHsPuokHDtG+2MwjuxaoqWyu3MeTj4lV3+0
omnlAhWqkwBMryPF2nwHrSVZ9JRqfZDe9TbJ5teLlA/+Tw+RXVrkcI+BHnvrA8Fs
42vMtwm+6Bw+2m/lGjuMRyE/5wMMiNxgWVww2bHkHxkthnY+pZfIlkzmIGqnpS34
40LtRgTk4N0N7n9bxrZO4F6II9zAf4rav4PSQpoAKci6SytfXfWa77aF5+ez8XUw
m6b+dZ6d1xkUSQclylxEcTTkkcvAViFphz4XHSmd8qLugdNqu6IU9C48FIU/Qf/j
NWcM78axKTDU8VVtCCy8cCDvMgbTm/Msgm2lWbWf45FVB3XBrmk7tUWNhEWb1Fr1
56LBfjLEFZajIhUiW2beZ4T8rrc1VyH3cwIqT1LJeDKa+rfr8/uOU+Wsea61G058
glLqIs9Wkksoxy/utI/3CUjbwT3qqATNI5Y9BUV58pwUb++9OOq/qAKa0qO12uhc
eu7uIoUf/BBbjyniCzYPq1ODyveuK3pWL/ymnZ63w9y4njiTAQq91Lx3r8w5cfWp
iz3tVrXs7nh6eRDEC0E0Pnm2TTcllyV+wlPx9+ChCB6Ha1HqlWiDVUkrwvEVUM9f
1lLlTb3JTpnAUHFpUdG1QAYpvrgpMtx27Q6sFtxvImE4bJkXHA+2zkXO6jWTNBSh
V5xpi4StToFrSXXU7gMQvcACGNwfaRQUT0RVyReexqV1iNMm7tcuWOaPjW0pUbYW
ar/QvdWfybn4WC6PGtUDq0uAa1ag4fH6QxsqNVsL0vSjXIZjxg9Sp1YD0K0lQC2G
82mga/NwcMLF5Zl3Rl4rB2GijwTvnBov5ThkC+lBsyEH9Zkq36qd9ZiwkqaSDs9f
KKf0/h0fNEBktozGXc+8yFKMyhFu6R+GZZz6LCKquyangSM32hKd83Al0mwwHkXl
58vQoq2qKNsb8vRdUMeRdyBd7F/UKyBfkKHgy9TnTastXeZWcSqhZ2ZQxxeOdDIM
ekKs9ihKsdD6e+Vtxj8dHfjWeagtGLINZjRYOyKlC8P9maydgrFNwHos3D0Ys833
hGP2pkBOal9nXkM15zc4GNN+PeeIjOBMQ42DiLLUBtvwxMXZ9eQBk4MR1X0boU+b
kPPxu7wM6czSXAzTcDKyADVaHA5NPPm/EbwUFLDFvWQ0rW5SvoNGNg7M6L5hc0v6
rWm1Ck2+LikN7caKiHAHFgIgUAVLhyCoCCiuiq8CZNo2zCD43KM3k+LLxEZ3jkA7
pE50yiLb4lYPi8LVndM0367o6S7sFKWWwH7DQ/hW5+OlFuXFgLom9IP2zEN/pv5M
wErr4WORuMz95KERRA6XTIz3uMUpEtRn3/R7a7pzt2p7t0bBvuiCONjeDkLBsaLs
dTdGm1rtEK20xGzsk90JjAEjJiiuOtufU3d66cccASlVoO1LiRgvlm65ys2r9bn1
fMGgzEWRl4Bek4vS0VHZogG+lG7H/V88KWIiA1MqBnckmj7dLdzI7VcKx2ZCaEOD
+PQN04TzFKtbnUI5nPrthsrYlxG2yQSMZ48h38QKMkl/AeH4TCfIW3HxGf9nAcra
gVpx35N3PgXPVR6JAdet7MCg4EaXkOOLnqe1zv9g8/KHBwT9xA1Qt9R51fYkWOl4
IEXJ2vUelZjTEXsuU6uZ4rzgS6xKSHMdJsLT9Zijm4YTHrwE6qiIgqdugvjUNp55
iHvaGkWALxeaOc6Z14qZK67egC2ZrFIhm/uXDUltHmy9v+8iPjqxvDYLnP8Ogd5+
0FbSDyfspsmUGiJuJUVHC/2xsnBBREM2HzJ4CIVb/5W0binx+/nbIxhTvdhnNGZI
mk7AxDylJwAr6R7DS5pXuBBaraA8H3vIntHmOz2ASvq8sMtajIFI+mysLhxrK8zA
rSvyF90luB83lqaqEa8CggxdHFm60E2F8xwnXj94HUk/xstgOYqhEVFEjaDOU5uJ
pfv4Gep6cB3QZgnoWF5i5RY2EA+a46QpaP99Cru9mIiOP0ee1KxgIZhV6bzrBqr7
pgp3PqdyBipaXEHiT9im/oFpEDgBwVcG3MnkFfHQeLY9WRwMuEwU4xBtvEGSWlkG
MI+8/p+slRtC4YuZEJbFwOTbfr3n39W3aBEYvX7MrQhknpB82H72UY0oUAC8PePG
37RILmaXsyjP36l4hxW11Fsaca4SQ3Ravg/wpFp9p/StVXAsXYqN72StZ1bqtLGe
xmBDRj08nCc8Zu1k/5ST+oHIo6R2Qj0sIkt1y2ZvD97DoFKWkuCWh3GBWnKLgmoF
r7YCxpTYe6yn+nkV5LbPxdwrB7a0wmyJnkY8woRLrUaaWGIEwGg2oSlqpsAp9am7
R0kOj9BEqDuhfGNI1dxmlBAu2Oi1z1KnJxH1oIW6FabKSTdLICdVqaFIet+Ic4qr
83kqw1LspZEnIK54lm75epJpZFnJCJD4qLhgXoFM5VXuzld8BBi5T5F6hm3Ev/KK
hoBlESj/ZM420U+VaB2wJUKbyZWRfK7HAxtX/vHgEmoqw6t288ZFxQ5WtCsrZbdX
Bt/Hp3a2VXIeRePJhpFhqCkyTPJMvV/swfYkeHYr8c4bQuI0zjh1xiSyJ4olZH11
d6cjdAAghcIP/nyMjAYiYPWMqdK/yWXxTK/GgY217/TfMibdfm+dIMppPvq35Pfx
e1GGIXM2ZBtfGbFhezXhe771VQL1mOGWbRswNvMmn2uHEh1ON+PX6ZdLiaXlgl1b
w5uEiSrqsOGtQWfa0JoJwdpUBJdZBjZipaTB9VeRE7DoJr8/+lq8Xjbb9WC3P8wr
s/2NOFT0wzirl9sw91ePyfF+p2Q2sOdknVgGT/7UMYH02Aqs5tZe3Tdo9JYSKgep
GwwfzS8Ziby8bFYNkbiD0afz5F18kJSEq+tFHTFVa8+5ie6kBY33LkiaKJZYJtsr
S6GK49ScmOdRmHK9Th//02W7QnTKMIYuoOqUgipRqL0Ts0MWzPcz/9STnHz8d80f
QC8kKSqyBTpFdR5O3SZNc7NSP9abfbwqQ31rZXYtnFBVZJc3bTO9T8aLYtgJ1jku
tdjZSqWg6UxMKwcE650w2fMGABQGIoCQYwYvaK01v3emsduBS96HJqfwonQh7Pnx
0FhK+XSgQ81zDRwJJ9JW39/hBoQCJJxWKJ7txMDLFzBLzCp6G1RPI6vFPxR/NMNu
LvpBgmLh+Zg4QurAt+vhFBKHxI1Ufqyf5N9RaKY+6OYvGjGxjCB9u8wZkHFYUuVN
82Kq2XFbWuPbd/xlRCeoaljxrtZuN5p1CK25AJGrU/mYfh+2ogXLX1pXJ+z4HQak
ZpXSQLOSIcrMy+T398RQzVo2QsGFYkkwuU+JWKRO9SvyoxNhjlnOVmqoUYH7L8JR
+PCPQVMqnbakWER5CxKbLEr1k6vnEGW5TAvE7KSp1zyWW4KMf43a+tkTjM6jGAzY
qM7UCtfaVL+K72YGh+6NyWpcwpxlcLzsCTjm0g98LnSckMzT2k2sl5o4+GnmbK+S
Fbj/9DYfw25Vcd/qPKAl4KdOrOeV8/kXhZ7K4Fw4UKpElQ9rb4x2AoWA2wTTLn3P
3z6naOCY0AgZf4gCaAnyUZsgjvbgQ3khE/xLAsmBtY1Lgs95Q7JNrluHudonun0t
B1RhNFA0Zc9wo87jSADAx5/h+RSoNF/huXHDfAo6M+nZfYuQCIlBljw0Jo8Dmo3k
A9NeNn19X3RBCQwaUIy0ITBwz9GVAi0U/k9T8l76YloITikbP/38VemJMRIymBe+
79ugFxF5I+s0qlVZrsRXOPAe24Y6FyDVsH00pspvX/+gAgWizmF8EDT0feciltCI
8Zb3w4gIhCq34tdlhRKWmAg8apfu4t0MwlUhg81TRJRWpt0L1FzwT35ZuVV4M8xb
VvmMQV8QYheV6BxJamVjfKkJ5Np2Bu1FAkty876raHtJSobHTPO0TgSHr6RMddA+
cr8AVTCRUR3em6eLFC4MuDw4LYNR/z77eUIF+Rt3bWUDPwQGtUwlrU6zj5YpWPuM
8F7rbV1RJ+shwMqTaobXuMLJ7wrKbNuHcnQxExxcEd55duh+0vS2taoEglMgWQVC
B5a5SS/bb6aYLdEh/lj/pTKsBNkjulbDiPO4jPP+Eru/NBg1UXrAcXa9zGHh5xVv
V9ki87pBQJZCOkgNrfrCUcjVnkyuilygWEEgeDPQG7M9N+ijl+Ssi3QlbcI962aQ
BhiDdpv+yewSt30adh+Cpf09ZbNBfUYwzRbXxiyLBDVl8J6p3Qt9+y6+PfWmIIz3
w9bzy1Wlz7hTyNk9QTd5abNCEqKWXYMzk16Kt2tIzl1GjgTnRSdxoXNUnxO75U1q
G+g5qZhc87ItLdRw/RUDSd3E3SwDvBcHHWaYlZoE/496EYK7wAlBRH+0cx36gbv1
Dy/7nBGH/jyS5d4FR3I/s0Thy0TJ/qAT7Qs16kTtbuV1Aa2foCLyG4CKsT/YjjmV
CCEArRZMgrG/RHNtu1ZONKxbOqAd6VsiClTl1oV5uBZe2f/78DkPTIsi0J58VlJM
W9r44PekahV+CfjO85AFvnVjO+77d3eVdMzAupD/4HRjehO2U1KmSL9ezL1M7vAH
G3fgdWK+qzXLSUP0o/wNP5o0WHqamLKdzlT6Qw5LsxVomywfKcZwIBOPd2uQPlq8
CPPIfOyvIihw6dyrP9kfZfXk+SrzLulC6pv0SJvP7KjWV78EUTZphHb6YTVoTLON
1O/GjY9bLZhmHSC0gXHcAT8spwhKR+L85VU+8JGwOFrJt9Hi4ip8hC8S6NW7n6nt
W0lUh49jsKFM55isPqBAL+f/yBhxZAp35v53YCnOGOOyVlKclBFdP/jlKfa5aEcs
UyrDDGiPIAXQteYwYgxcdbYRUZ7AkfmpvM3VJuPI6mKEJcKB8YDNaLXVOsyFJPsc
mHcL2nlfhpZhcWLJRX4y6g/kW2UE9Z/O3l1y+Il4N3ubN2V97TlC3K1plyGJxApM
9lTVK3zLtqXGI1wmcHPGHjlQ7OHNhCm7iBAvk5iUtq9Kvh7bm5mNN2C+aiUOqJFT
5gxr+uTCMn+dJJLp3FgQjkDSREjscXZ2CDdrmnmyoYzaK4/0fRrzGAELXPPfqKX6
i7dYgZ6ptSz1zlD728BigTenunXeSRNfgmG/Vto8dQSI2sm6g7A8K3vto0mU4cE5
73TgjAXtLWgIfne2Oy5Vwh5uiTPpgScHMX64O97MMC6jomgrs48SRM8YksuhnFpM
YJUKNNnxxcoc05w2H183fzkAUON5O+iIRgzEp7Kr1EHgV3y5DxaOVCRB3+DCzWby
oI+gmVtKvPBqSCtEqwsXQQBCBep06wLpMp5LowgjTYHUeoAQxvxRoRfC9RH28iiY
Kp39l7omCuEnS8UNFOcQMFhLQWUrCLiKMquoTUZNV6dWR9Td0rp7nbtcqno7dYZq
MnXpQfX0+0zpPWfZP92ZJi/RvHNNfiBnEPru3mAxDukqdTeWyR1qLA6tkEkxsU3q
9RndTcIfU5/asxjYwKpDL4+ISWzVyEzQYiFvAy9JyEwLxt/mkNi53zRn/4GxNxqF
Ehvl2qAStwZZvFhpjEMwXU0AJBs38aERSow1u+gXj4U7aau+izLZ0OWqs4iSleGo
tJWTlkxt+E0dxh1UQi2TaiHbh8YRAcdZjwyaIYwkkizGha2RBMGXXlVW668JRUsf
48xsX1ISEE21FMI40so5MtImqef35PDvt/a5WI1d3SbwXlFvW2npg0xix5AwP2V0
8xNYz8YRsSLQI66UFcGZ+dez4ThzwJhQ06tZ8iVfG99Unv0duUm6tLkPlAbGNlUh
liW+If8jGBZ/6mfbCtqdJABPmSbBFE1CdkDheeK0Y/nXXRRzL8BOCqlGQtJerZr0
rfCbw93cvZmZ4VJ7843vDzP/b9y3hLE9V/Mz0J1HfD2Wf86SqvrjcvP7hRc+tY4K
GMQLiGNpIEcaM0JJBU1rRBeMiPH7MDbAr+kh0NHvqyQCBQK5vEk82eBUY/wfj3Hw
/acNTaDMiOnnqEIOVExgtO4OsLZGvWVt567vCuzEc/8FNDpMTA1YFsJHrUmY7PJd
i27Bsc0ofnDi2ylKkvuaxLsBk+CcJDCilhniInUgueVy3lStZhcY7qQBdTOLCYL4
BaVnjABKS9HttHsxweLXBpWkMmuAyeRoQXMSSrYLWuRcIb8Tca61og14y5OPl7XZ
u5KnQHdsyXm7pAovDeuh5u3c4+Euak3oSodo9KgwpXaHN2c/YrJa1p7ZLzE7GPol
Ablom22eusF4KIoGVj9HnGW7NDRHQnmDI9aPVIYPw+1xQfbG3bDnZjfNxZQz1+85
4O5c+7E3swV8UJz69HMkR6WLZwaNk/S+eNyZh8wQpqntFaGbzu9az56qsyxbIA6o
QtqKF7awsQRoP1D9K0oSwtRc4RJi31MF8Oyr7yBBDeU0b2FJGwRxBVSgX1aC4WF1
vmjLC+Z9ZYK8rdYU+MuJv7Aj2KE/vJNLW9Yj/vkEAJPQfYpCS2UNQvn0HVwNoC42
9sc5kf9M87295QA0Pc0OdUEsBp2FDiHzZF/FylkeMS/+YdRBmOMrLaHQ+pcRXKOr
/rrIINNv31oJuDEmelp8IoOo+tGnzVVMDmAAeiV3kch9eHD+Xq59Gj3gVocwHAXC
COsj9KanAQaT6S+hAK4PiygAi1eFFstznqsY2lKQBRsgkSGKdhoI5loUHsLQZwMH
Rglj1Ieq9e79IWZ8QMFpI8fW2A8VrSOfVgPym60Jk3l6DUP0Z6MrxC37K3JNqxpu
YQWYiRgK7lLawBbpym541xFjyfZtba8DoIZmU05VrxNrr/15olLXc5SNuXqr/dpw
wLEsLCAAf0yYbu3psfW6CB7HPqP9DfsyJPSuDgikVlhVYGntTgbOr3tbuQVgNPlJ
FG97hK2vCFtqMKO62zVbsT7NZfgdrLu6uetjL+9dzC/iJOItBez1a2NCPOFy7O0Q
ba0kzwf1aY9xrJcLiBZcY/VIbrz0TKGzNuv2AMpfC44humi38OErEx7DbWEqfuNE
HuADpnD5uxxNPYJvmcR3/eHrBxPBKqZFINOwRUy45APYaaxdxTXS8ucJ7JFDG2GN
TbeZLOKA8iSzn4rKNQAMyvW1CoA7aevkXpS82Y3a5FKMX89XhABgeihTI+0OzCYd
Tz+HTEqZmiLzuvgniuUyxkUy/MfnXn/7W4pB8ufDRFHO2OVynEc+2hvV02cYiyw3
MVO1WAz/TP+SUcSvCK8AGJiY+nrPr984AeATyPqKhAn2ocdrkDOwLfoDr6l8TXt6
0gKpBu65iYEnc3CqNfxg31x0aZypL4DY/weGCNHfNIxWzg5KsHk5L/XJDhxYxe5R
ZRukgMdzL20gfpPBqsjtX/WSk7qYZfG9rVXvTUlDlS2HG20Z68pMG9e+Mg8p1IZ/
VmIFz79EcUBO+VnWKf5zdHPRm4CAHEany8KMXuAvmk3HRnbSk4zL0j9qnHmgEKcu
J6rBo/6/wGWpwUnwMk+qbw3AKhza2OnY36GEHJC2X/qyELXEmZxBhwMLJViY5HdT
UIHfnyz+pWfStMMLKHmCznYCC1pWyXn9qPFtyj5H9V8ZHLpvViS0U58fYr2F7eFa
UCLiv0eSJXghOP3MkLVbHbbyPlJDgBr9GxebgqGhdRknw/KqHxmNhMXSPzlciq7D
VHcC4dSkZCYcoPIMX9juByt9fQOo2SeAehf0/GhSmqNU0rMejfaVbLlroHeuTcN3
TuKJqSz1zZsNhEr/OAxibwKywyo8E+Dve4ykAGYEt21et8fmD0iq/mKiB3dTMJ5g
4EeSQH9QKZ1BcHr5S045Gqbqz/LkHPbCX3yKIR3FR1F0qwnchTaPms0hQyQ//JEJ
/8EdaA91fPB8sr0++sRmImIA/dZf8r9uzuo/8oP4vBmcmd9OdrVSwTPyJBwU9+dz
bL8RlQ/k7BdkBvi4P+JkdQo86hxTxC+fjAwWwKmkNe2vE87z/YXPxKaU/IJ89SQ2
rzaW2feq5afCv6CkhyO1rwVO0FypCeaPYu0kG17hyuwcRhGUBjBe6Rax8tdO6ZP+
99/Bmah9nKs8tAB9mWmUkWsb7wU7wNw620uEDLR0T2UoATVM1mJFDlhXNAnkSEnk
0Y1BMZBinPu+MeaKTIjqG6PH2R8ABObmmE1iyz+hxtoiLrQEEskBDozYpCX2Pqal
wH0LwxqkvZ/Pi4Oadb1hbO8jhKGihuCO5WVDP6kfTDExsEcpsTs6k9ezPEr2IzWj
/6yNz3ctByfJdr+MQA3F4jV1i8VgWe+GBWnH6RlT6gHFH8wv5xfpJMLoxWU4ya7S
/ziCLI/SZTuRDNyI7VQtojtUKyhoEs01nsUN/e3EgifSVE+alCjFBkX0wObsgnVq
RnY2idF7KRoH/gT69KpxeSzi8iOfsK1AYCQA8zj26bDIDTa26pH1El7Qqf0e/2+D
9d56IqLPgIN9z514HuszBEcjxJP3dudjkOpuFssKebUt+vvhoz+ppodZ2PSqc7MN
0OU06VNoFSVGxHiP1/KWV2B7WpQqmTKioKLIBqIxai3+z3i56Rlc8uH6/geNFnKM
W/h2d+qoD0oYv3yQ35Oqgdmn39d6udGRuIuOgq7PQvks76KlAuB7EGNTZJ6DEBZE
Ene9L+iIuw3zZaW/gTyGAbBjVjM00+BmMem4mXPURYiq15WLK4dWjb9zyc685Zes
1uavB+2rylVT9KeFVxYMh7M7y9PFoXI6tNoDyB+n1RmX9CRGi3vzct/31uS97vfM
U+oRR0LjSfv5qeX/n+LgjDIPXRVrNSXNbsPd2MiCih70ZltB6RQom6k9UfuR+kK7
Y/luBxPJh28atFyycrpOCH1MXyRRysS1heMB+IinhMcuh14cn8iUKBWh7pGzIlfK
LseYRdU4NTT5Tw0dSk+wqJ2zMZbILXBQjzbRlQ37y5VmlYuELfZvHZ2+aQGdLcMk
kUKNF/f2p93oKdRH1c16NxcG1Ear58x0GobF/zmAP/VsnF+soQNINKIbBNQs97ty
pzu2N73el4PDpXYftvp0yhY8z1zMS2QOc7iZJHgkWpwH6aGWUaTgr3Rq7H7DkdF+
kCs9wmyNmEkqroemoGlw4wNBKCEcuM6FApWpLV4W5v3d8oUmoKHAvIP90EaM/DHz
8UNI2l3T+vYuDZ8q9SmpGQUk2KWhk3kwxyNayBSxvAIDxypHyOJcMiNdwqPYxe9+
Ase5Ev6yw3tHmfVzm+a63+VlfwF7xqfEOLsVytW79IIKbHF2t3OWeJChskXRk6W0
ARaTEY7MQiWeRov8kGMOPsdb6Lk3B1dJrxE6MQlssDw=
`protect END_PROTECTED
