`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
s+uFV2/LIKd6bYl3CZQh7p1VmwUs370ifSSZl5Bztm5EUoVK3iPY8a82AQ/bqHRv
G4BUKMiunvoNQtYA+mW1/rs1DrinzEMb1J3eHTWIh/gDSkvfQIPFYENk14Cq1+rl
/Pj0+4Hd/bd66GtrHc/Sj77ZHT7tCZqpIk/lFU/SBg9kNdM4MJSZseSOnU3czN6T
wqtFa8GQa5BZUO+opUaYPjjm94Z3XCVmZQObgnRan/wSGykr5WaynVm7gmP8w5l5
d1kHwNsB7B7jdnTSQAbvYpAm4EhmhtKtOxaKDmL7HrDJd0CZJLEmOqX+CzU1U6+c
W1vTZDIoFFUF8haXeIQLxiUHIyYczo3MKFsyXgWdd0z10yMHBGeUPk55gX5AAdcd
0ZHQiWb/89a74Lpd/Zl9XX2s8RDunAFDH6vJyyHGT8fUTiRlgmpWw80croEKnYTE
yAdB4dvPitWmf+tP2GwAKNDzldCKe8TwqlUlGRLh+PVGvz5bqk/RssKyFZSiW4MK
oGDFXK6zQoPbXdc5FxjAYPOzrqpBY5ie1cMDAtfhAFDG+c23YDWxTYRtzRHTTVqi
QTnsw7H04ryUCQWgnnt/Uh/CdgD2z2y9i2edH9ql/0hvuQmwizVS/i3vRqtIYh0b
H4CM3qhOExE39pEdVUWKVaLC8/LUMaS+dqWyChjnH1vRQ8Lw4Cd1lltcBY0ydL38
Z5h+GKFsbsvQ6LNaMNkKaT27j+++qT44G02FG6ZLDsfXASGiRjxRfa1LsKg4rMLn
E79xH35xxsOg2aliHzQZuEmgMoHpNj9gV/2XrWG/8haoJk6eNyDuYdIGabgOuTKZ
RwE/PkchsddBQVyBA7YmCEcDuAtiO9kxU39ulA5YqLEIcnv3mKFCHU3AV6vil9iM
Doeb6IM05XI2J4h4viAMVLRnppiNcNr5+ytAa8yxr9oWY9w8hqOv73MZSj0XBjqB
ZBPXCx8r/uz0UomAlkmDCurpr7RQ+fzVR2iP2jOR5wBuToDK+glg6FwJnPCsl4uv
6EV6OM4uWsFljqOXPvRo8PuV/YTyJCmj3r8aXmQ7Lt9Et8NPmBEh8MdJVOUsnciM
9M6YGQzT0PcJOZmLbd0VLmRhcoybSPvSRIjDrBG7u/IsQDJTZ2NZ0Zy5s+/YwJtr
hNl739AfQtAIKGLna6oazjJXIxoi2JRkxv9BXVrFXzxO7DBz3ERdflYG40C5v+y5
vU4S7gzHm5iEulEsu5cVi184jxCG2IYK5E3L+Uq2gJHsUrf+SEnF04X3ol5Opnf8
PohowOs1hiuYfls/XgA7uCmAoCBA4mqAuNoGp0xUduEibPVUsXz51wmOVG9iGW0U
MVcFPL1VyqmkMbYCvIx9ahxnAXN2W/DTfUerlbhyajjV3HJxtJTVQg2qfv0c9Cmp
5A+XmPGlnsJjf98sRid9rUT+HUTmnIfOo21hghgw5GKXMEeZwkUxSa/3i8aXuKBf
gNqP3NukImmFHZj0MbglN2/NbJGNXYs4hdIUfF7dKn7C5X/Wr2GOyxuj3NayhcLA
ao919UpPGJuCYABs/LvwsqO6oepuVNA55zzcWVI09rwqyiucghKH8RV4my3laEKr
Ia9HnZymI8Pn92gGdtq37od3CPI4U38hTQJ52y8dKFLcgzbH69vEj+ZiSqHFVDq9
9QMbsXfMEl2EL9Qd72O5VL87xLbAtUUCKUlz5yyIWQeIJpWfmk87b4PeEDSAJGmF
rECCaEldy1fZhcAinxKDeN0LuCk1XhZ0as3Iiu0eVQk2dItyeiFWh417b6MWORuv
a4Kyr8XS8sE3oaTi2tKGynm/x+Zpldul252w+0ixnM+lVFrfqK9tjKgM0kty0HP0
LB0xiEuvHyDtuCCP9a/4AuBS8naBrBKDVKWB6hbkpo5uBN8Y+VDqzCeK1qELgiy5
sruby2vcWag+vOG55dmql6o10BuHxpFu5akbgjtPQSwOXpJtyiPi3NXpTaJ3LUsD
15zlBbRJPhCsS6r95yqAJ4pn4HhcSMbIA41zM3J0f/I4g8gp4xNYMvot/NUmSdwy
FX4epIROWkrJ60WdasEGeDNJTkhpIZspEvEux/yfBvcVwpXQs6HaP3zXT6fPqTUN
SnGQd1tj/XvWpGib5MrAYFXzCXJ3BiGxt7akLJcCoeKHPRHAKNC8x0AG++5ETRl8
9WFQuJYhBMjMOyXjdX2cX0I3EM6qSyDXE4E3220m1Ak/scqD4vMXXKBVqRtgD0qw
HG3QdRxd7pcXE3FE12+NCQ==
`protect END_PROTECTED
