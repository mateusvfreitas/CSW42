`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hnhfu7ePjcNUIPJsocFRJH92gBifpzNlddLSK9NTdpMzA+FtJVrq6Up0RNVo+AwI
e689trDYvahJ77V/VVcjRT8kUGM4P/5rfr3bJTR5gFCKpuXefdCHDHhZ1oWA8A0V
d3YiODFmKGl6jgKrQdrXE4V5v90LPp7X2AXPcJ6oBqCEArmOOGJsHGutArFnJICF
f54s5QIh1SjHuUNT5IwbxmOZwUoNeMFUkFPL666VKdGbislCmJst5G9akdRrzGbd
Vda1ddRfS8Etg2zQpRWRWTo2vGScK1NDJPlRzxZzH0JhVcduaOHgQqfVDMsVZFyR
2P5aA0+7Oy1w+qGf70UZb3kxWRR6/UWkDwpEWijVuFI6zug+T8kstTTfF7nHQHla
+/KLE6puFj2IhtE0cDyLdbPFlcEv9qgEDGPcsOVD+/vflFmNKSWZL2ek9R4CXJO9
X28Bc1Iyr82fCUF3FU8eOrxXUv+geAOOs2/Hqg44SmQuk8eOFkRbReUfd0kInP6k
fM39THcYM7sgmIXBL6EoFL+AIZiGziso6mZ4zWNoort62i47AvH2yDoN9qs7ewTY
QfohdZDMzeNt4QuwZcq5rFJ2T0lcIUXBAvgr6q6Z/sOitWVTBSbZFknOtDI6o7rx
N7Ixg/xHTHYK4vf0fzbEZgQ8rxLxalVmkVnyD/0ZewESQSr0R3sNGxCnAKDyyTkz
DHRYl+TPOFNlnr9RN5zhIbt+5gTYYPy75ijIWkdW1VOxlyvddntOFhE6pBnYodiw
RaP77tqint0HH7OmQG+qFPrINrD+K8s2EeGh1FD2wd9wuuqKMqvX9Saw4DjmjhFn
NyDWA+Lksj9Wvt8KIm+m8od2YHemvmJ4QhrJF29zjkp1MspxbAESnQ+Zobo1nYMN
F7oJ187Hrjv29lynmnx5UmNY64mgXoFAxcIhufhqUZZY9Ppa9iCgjmGB5Cv6QzdG
NBPsHzNX5auU85JIqWTCdnvQS+OZJlbvIkeBJ/DLE2pK8txsAFnjuqstT5x2wLGP
3aBoZ9+lIoyaKezw60+yE9AeYfvDNDQU4mjC7kLNpQfKXaw8AIEi8QyWbkDFT6gX
LRo/f/T2uprhBp5AJGskoTMucdfK3DLq49St0kpuKUKIXlFTKFImICXBgUACRR6c
Pikvrf12i/Mt0BmLhJC/JsSA2jL3CvAPZljszcXiqaPZTnybNxdbwta8MZ9ZTQ1h
ke0CVcFRuzV1obbWHcZNbXGKdfDd0/6SmktokLvefjtqdfyq/I8sCFp8+v/69iBw
mzrlPBM4S1UutA8RNjKEnKWuPcVxHyzy41Wub+PfvuaU5EMKeK1Zv78JIzlfbDst
q3irpmlxt1BcYibYZtE8SDQyHcAQiyP+94nnM7iNmEwJZ4evyfOKLq4BcxvY5Hh6
AIxm0+0PnLhw5vdYOWrOOEzzk5PWKp9BnG3uNrl66mvRis5/xlHpJxJv0ZS3rapG
Z6jqqpcy6oVwmTWFG3DhV9mgADGYlgA6pzJgDxKBed9iiujC1vRv0dAbr6SZNk+7
h+tbNj9ZWgeKvkuzqaIuNFDfYIpwS0iuxMgOn+3+zLx/KjxmfLaVi1SYwnno6Xid
2AvwfG8Yuv1mV8ocKpJUZVhb2ia6fEBU8raLj7rU9RiI2KCoNj/aU+nteoB9FqTt
3f74yHIePDyK2UWyTdxTSWsfJjw4dYaYALwIogZAzUO26U5quupGXQqzituxts29
weCu70uG7QY/H9aKOpzilMzojjra7qEsSEs7zcoy+Mwu0wiZb6p/C80DMzS8+CgK
l11UZSVpuNi7r6j2g+UAZIMA1Iz3L7wr5pX8CB/8ahCqvdVhqjZ0XtVuZuKrUjia
lBz1HEDHHU8qKCuMW11uEM24ohUZK6GY3ovHQy4zxvwzHY2n36XvpxWoZanOw8mJ
zO1SVeVxdvCnLzRj9FoOImAxdD2l9mRgrbz9tiIX5XBfjSPDz40b9SR1g7LLhTkE
o5+UGcSR3V+mToyhT2m2NFaP8qRVeSRyHPpPQ1IkrEBpg1ifSMyTv6XI9xrYn81H
EXxCBKR9dKafbvloMTRM7Ffoko2Y9egWYlpwCa7wLor053Zb7KGqZ/Tsa+15qx69
vgVLDMWAZsAJpB9xDra78CpTJWjBmITqeNqZmuEZTNZi2YKdD0I2biO0g/iiu8ZB
Gkbaqo46HPDkMLnuXTnqoLqA2uwRu138j1lhVCiUCB0xeDiMQF6kkxJWODoCMhTo
DO73GPiJTbET1ptJW5sFowffG25/p8d3AP/5s6kk3aCnglXxg3388qvlcF5MZ4/J
0ryUV36naGQ3YN02KKHmOES/ta+xlTSWFfYhM4hQ5Uk2Q1Y2/4c94HfwKOCqg76x
gQxEywIGufNk3fBdY0t/1sG48qxcdwV+b/n7oSnU++1KlhXAhLl7LsZoC4QxLqv9
y+/YKPTrcTDQ5pToBaQrCSYUV2JmTDHCEWeNLUk/RVQFFC0cccCZlumLpSJ3/2tq
n1lBEsMbyBDGpyaoJaWEAIxKCDBZWRShpzgL47R0Q4aPp50GPsDAtt52iipj1om4
MqPvvVOz0+VSrVrItCGtuPZaT62daz+4YaS78r4B6Vdm3neYtIIJdFaWCC2OtiwB
egrWfr7FEXPfXMIVdEGXf1mUByXguH4SzObd75VpDb+RqqSQR14o6aOfGPXkwcLX
/CYy7rNLALcnOr9H5vz7VysLuQAL14fivg+4QW4chOiUfEzKUs0FaemcROXjvDFX
LI9iIk2meLIfSJ8h7ckiLTUzSvK8yr18A9S7inq3oYujuP7mBs6p/W59Q20gpL+m
7iP8CmcAYPoV8JqiejSlOt0ok/W4miiv8RMsb1yT6aZkcLQcdkMDMB62zoAmvZvH
yXr7oxq9WfLubfVoY3eoPgmyGnbonmCBd242FB+NurAt+VR82Oyt6wmw3b7JWLnm
7MJG3ZUHf6BZ+iMbqzu3zQarmfse1nYlqT8zK7q+vDrE4Vw0jNxC73TiMgc86dp7
Xifly9G3JxH3EbSGExfMXf4mH9WDQQguhOBEdhh20mz/51w5ih4G+YSBbklYiiL7
9uXqEKc/rsYaj60/VEsOp1xCnxuoHnZIDDLXLuvuD9UQ0nVk4YQXDus0ZzxzRj2H
EEooFeR0FTMsn/9QiXoZ8noV57XB2wPOQjDZEwVuRmQwAuw58Yq1E8m6Q2G0nL5I
3FI5EAyYKU3h5614bZ/WZe71MGXQDQJtOrMdBVaUz2jrxvYVjtEFz9uMhJkaBRcs
Ms446eCZexzHg03p0E5pCUzTNtu6OPC9qshe4Uek25OQrgawBGQrPTh3s7i0VweH
CuVH/BVDeFJqtXU3S9baMXU7N9rOD4CcburlMWkl8FnMbWH3nOGMtJX17bPJ647J
HhvI84um3ZkOp57aOTTaeTH8LtwFvSqoB7GD5BO2WHbv/BSBUgyqJ99Z6A/ZE/bd
wvBRCxjjS3wMbLHVrl44QKINJePcUOilK4jvo3zolNa8WYgW5DYkltVXDMXne40Q
Q2tIpwb4Yfw7OyrQ3DfDrRKGqbWwBL8ZiT8hfEIDlrCsn7Gom2ZjB258vhJjoSrw
Uy4q1XaVGIiobGFl/clMkKkNnRGptHu4XEItVBJZzQdVCWMIVgbqyBgNFTDeBG3j
6rB51IE+ALBVQ1TkwxxkdRmyxiyqUROZpOomstq8Vf5k5jHnfVFvJ3j+jqtVP6y9
0V3P+F77evLPD93G10WBiBmmM2ZMIJFYkVxms425Rh7wvMwPiwj62WdGoCieqIHp
R2wMxSiTptLGso+3+PuSAvMwfJ0bViivPXQeUkrXX0507yKHKjQU8EG8ysqj/vth
0A9smZkLiQ1iOmP9dPyhYMUj02NDOM2aKMAlzYvqY/t+Nyi23qDgaRidMxBp/Mzi
rBPWIY0xnOGwajBu0Usbn/Zra9sLNVox4IZHStlay4FZCfBQBM9UV3K5nPNfk9Vh
VIuE41LXz8RRrP68Q5Knm8r7x9+hPtuTp4Sbiv6mOpZKEe+nCo03fUfejpM3mSas
AM9mu69UlmsIhAd5G5a+F407W0OT2DGfm5F12FCFKrI2kC9Zd19k72BOUBpoGwhF
k2uUijHV6x/hH6GuXZdXtIssDwoQbHj05WEnlBoA0CQZLeLBqY2J9/5gO47K20/U
pmmKozSCIslMog4TS/ZXFUEi7SlgGZPdXV2CM8DxIhrQu65wNYgdrH4LQY/tlWmj
PND8udyVhS6Bw8FejZU0Vvjfrzqsr05TumT1I8zVsG8ZKlINhFUun0GvGYqPlzYZ
8PUxfDbEUy/3/+XoZdcfq8Ln1VoQaFphYLwW6vBXIyzuNXDH2eWniEjHzZoz5fYA
Z3L+IMzEu49jg2Iw5XZlgMsY5jzXy0igmUPC9kCxflY3Zxhdfc+xvMju5x88vvL8
eeFIr6FTLglJIobeOfyKGomyHosXMmh1SD13msx5UYxkKF9D7pRgNRsmYMAjEIma
X0HONyQsERtlOIh5wkFNIS7S/9aIDi0FL3JO8Crgs8+wdf5YEGDRcujuPSuJmGWq
eY2liL/jjTh2OovffvHzragYy+DQ+K1gTDBAQ109zUSYQOpTrMhNzhVNRo/I6Q9M
opzp8lBTUct7OF/H+ko/KE4Q56/fo1u9wKZTlJbR193ItyqI65DfxE7MF/pl0IsT
sJQyPiDOLL5j48Y6vUPRp6uIUZT59MSo8+vftrcmG359Ii+jKagKiTQMZ+6vkDih
CX9+8sb9xbeS7L8JbAVbJ/oMx/4tA+JHHv+qB6a+edM+ab3ADepajkddJjLzKX4C
Q177t1XQRwWUfzAJ+9omuwVzOrCV4nIxr2HZflXMoAy4fBSnZBVQrJZQ9vFCLvXW
5pgMDfDA91JJZHjnbDiIsdedmX1x921/WlqCEbpQGU6Cs7GObNwXnkt4Vlc8Og2u
SkdBIvUgckjateRFhtVQjYam1TleMZCLNP8KyqLQGeBhrI+13SPhRMcqjJdQ5GC8
TKU914ZuLLC8AT9LZ/iF2HhsuxxOC2/KYLrBXDgkIqcWNFrPDAAYl/eIFU+Popom
oOw3RADZ2or6wItJ/66TCbQEsSsKACf5UqB07kevIT9zQ7C4KfALwTYTTLf6OhNx
vbZoSyGcqvIdEh84RtWE5L/gfdOODfg7je2+STut1xg7NRWfB/s7iWq9bGCh6kaN
ju8oC881w0w6a2eU5i6UCtAv9ebnouQ03lsI0ANLVzQxyzJzq4fcfJ2E2drqV+Vg
qas9OvaGnk2oHs3+Y/fYOcEBbS4udMh638BpxZen6fSLCpDju/tveZ5IC8cGaEa8
Gkdl3+EWZ1ru/JhOxoV+p9hRSmf9ZiCnOa7bJxixVpUOdRR9N78giX4akOK/WpTE
HU7HGnVmWY41R9ux7TD6DfQEHwx3Zg3UeZUiWzWTZcjAcamm/WCeZyD5TT7qcrnm
fYDZyX5AhidQ8380LmFR6arqtCW8MLVLAtcB8p59xg9RZUg/632u6UEr/qdblREb
oul8YezBvAYsaMiqdWqegOYT6Nt2S7J2Crd+QztW3EHym6P3FNFwB54A5BgApQz4
tgzGiqG9t/KBOAr1O6SNRCbJJrhmfU9BWTPML1t8gFHX0HGlI6h5gmFP84/cj/QB
n2ekAxq33on6rfS42qRtsalOP0Rz8IV6NWiK+qEt8J5MzL4A8+HiOMgmi0H2lS1r
bIUaTBLIvRHtuBnXJ6xGY5IX4GxZFImiJc2a4c3nm3kU1fFigSz8t6h/4h1xo3e0
z5u8s5J7OidO+2daVajcuTs0Fsp1s5Yk9ImQDMMskpYh7I7P0rXZE0LwDOfP/LYI
kd3n/76DdRk708OMQ4S2eiJ72ab0lLy/vM9srAzQMK144kufl6BFVTr9XdkQ8LUu
ISh4ABz34rkoY0y+Mj+u0p799gjmtOjVDPlTA55gseoZuBXVtxxtAwG0fYSdxjrG
RA3pUXgYGMy2J3tG0jKI7LSwPoulv05XQ7vbwbPndY6YX7nNhIDKHyTX7w0s2DAG
+26XYCreWyD8MYsH8WLjnZa3OQJ9Op/O+jb5zmIg9ulo7l6oxbF4+ivD1mKlhl8I
QDldQvbp5B2EZgpA+pV3mMVMmpbAJOgaM7L7LSd4YovExzixYtKj6CqdXHYfmEwl
32oEQN+/FwW9qiTI4r8KZb2T0YkIOHS/2nwYe2+5Wyry976ByoJgLjewfbNsZM/z
BQFZENbfpU9xudG8kjczdzrBtL9D6/+R1zVqnvkw29EJGOJgfVMpys5E3jzpaaJP
8yMaturHldgv30TwoiGZmqYlnrYiRynIAVslwbi7MU5XhlOAhpO65IpBCx4cM71w
hBw1tKWWbVOcCL+TBk1IKymmvMVMafog93qebyrw2EecDJLUNUM7OaS4pjBpnAP1
BcAAZWsjnbab7z8Hh0IrBoo5P06YihcrSdbB9rLmRymNSZ6iZ6njmzp5vGBbWLvZ
F+W4ZbLKHFhoJOdeUyzdFZWcg2QEHzSW0rC5siWeDQ4hczxZdpaVP59tDNsY5DpX
SXRRvh10N/Yzf5ONXZYgTLRMg1z6rHFeQ/3FrPOxgn3DPWrEyDimG35KzsvQxjAb
g3imOLuIsmN/L1xNuRGTaznSN9lXwoWJg4Z7Rcj7DDpAllx7iuedfIZAa8oWHPMc
Y+C56y9P9nFEtzOXmSCaqFPUOUyF8Ut4yPGB33re+mfMcf2h+u+/B9pM5dp3ZGqn
Jo3w+OGQo1MKw/Jd6gDNZfzuJbfCPQ+IG7eYGZwbosyZ4crHtpUoxVicFb9Fqqzt
AjTOeLxtGSlFwqa9EfifN9Z8kTZ4+i8nWaYYJQ+dcIAZU+aeLOb2oJH9g/1fSMDZ
jNRIzz8PVnbV5AOQMZ9wGJ2vIulnVNqrfCuZOq8SE7wuUK0NUlSRpfgJO8s0msyG
e6mcj/VMXTWZOvbnAK5yeEU+sfxsPHaOuV2EWsUhcOcbGgV7+JdfeifMF3qxQ/4s
pByl8AyJtgNLpInWi1QjOWYO5hxABDUONE3xIsgN4qYmuAptBvufosFOSRi86fDe
gbPVTo1pA3i4jQWRIa8LAoCI/k3coQeXCx9fOACpRb+CFQL7zgxFyW3hKovmUsEP
FaaNUJ7P3sChm1jqLSkpmYvSpFi5UkjYDX8CJQg5bmR2L7gB7pe9nQjGqcD/JU6x
oXNtLgMFvCLMwPiEV3TtKiE2bK54OMFHEqcXHw2laq7nc8n7AjCYbSk5YqrJXwEY
B+dfoQIk6u38qxz4E5hM+m+9GfEfQMEubZT1PedtsMWQtR5W1yw1uta+laK8FTd+
zCSij1vksrwo/WXS91ZJThXmhqpntCuIpB3TWQe7svPWVKDWpqkM2v8Br0aCxQMd
rhdbNL+vt8MhRH7/ydtCg4cRFYav3cOsZJo33PpSM6gb7GHxSqSNYWaNaLYbqWH+
gYVpKxGC17z6/9xstuMN1vR+h48H+H8AWwnN/Xs0ZXtL9Q5H6i9U+t2+/RAdnmZx
pRDSIYQvndjieko0zhucmVgOFhD3sVoWthmEo/FjNTNm7uaXXZdCTzMnAm9eJnol
YlNQcndEGZ+lTfhdQI2Ebkbp7vzDI3eBPqLe8rkohgPTfi6dAWP3DaAgEEeASaJc
db9p98eNbmPfDqUmFmjmgBOFUei5esUx+3ybuOBvW75EE+jrCXX+QfulfFaO3cGk
J20C1YylZYLZJVdVy142KnDtxwoeaMYZ9+T9oEza8BH47B7YCyYsqL8v/Do0ICOb
R/RtFXRxlydWwwjU/7lL00+R9bO9O5PSbTcwwj+tglbPJCgY/K7ER5cbkBWSS+Tp
YHLWK9ShssuUUWBflWkP/BlFcIp/1VxiQQDSmUFvT4d1Qj1XgYNlbvyjurmQZul2
QpWS/6eulIj+m3D2UtwGa9S66JtCWokHany6WuTZKUFrHwynrZAnCE1zv2O37AgL
0wmtM+X7XzL4NpnWMwo5mg59Dj6S4Nm74FIHmycgIMuNNe4tMQTKa+QJZ5YAks8J
wv4gE/QYiesTyorJgqizbvHkPKfHKQIfGx4hkbB343VdkcI5mSQZf9utO/cyMZoH
w7MIJDCMCkb9M1KW4av49OF406HPxfTRj/yRb8uCtnYheGvoEzZ2t7UFjXzw+c7g
rYcJZ+52Vep3IvoR0zKLBTGix3KJErZB2SuxUSQ7fxvy5w5x/Mm6ICQzRn9pItlr
88neXkLrT3vVvRL74JbqWydZ/StfvjqLMX3YIangmEs0vhaUvZZnXALZNFb+uYGq
XRkocdUHCHWAwz5PJ5Hmfngz1H/IoXbacLpdjTBOR/VvCTzbN0tE5s3XwwnZ9mtW
ul7S+pOhspY3quLo6q4EZ/cQrzMVR9xGQDrlI3y63UKwqdRRE6JET5HZiJAIg0xn
rpToXb8r6cx3A3+JTaCuT6r+unaIG/OHDtQO8wPQsfH5IV7h9/99Mx13Qb+hWgvl
gyUJBBxiTMHUW5ZstuOnphr8buyKHq75wQx8JcZ+OLh/LVedlaHjBrsG0DzYzEgp
1XiqueyvE1lDBwTOUQDk8/7s7nxc0/2TkGKF7LWcM2CpnqQUQZ2EwnwqizTBKS2c
fE185Vnxkt8Mn2o1TltmZhPi6Y8C6sKxeKIixeSWYbpKNvn8gric7VujJ4XndgFy
AGmZR9NdGT2vVAh75/46NjyjnHZDtQcY/f2bZqW6kAz67mNnq0Fawp6KgUWgLKY/
sNeGcv2NcXbH99em9agMAvHm4N7G05iKUzcWEt8KdGfLU6eh2/WnIrPiMt9nISmE
6/XmIYnrhu0uSb7zvOfTiqVYdT4nj138NEX1BmiadwJfJnIyQ+GsBCZxUNumKq4u
uz5we2V0Xqv8wolROrtw/zE75UJY1NOdrXUYz36fIA+OlmI68dKFXDaaABRJoiug
t4Lu1EsswYZTmPy/Oj9h+D5V2zjYuFV8eXq5Tz6GWJ0=
`protect END_PROTECTED
