`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
gmfBWAHlGP0+0MIIJt7q4W+sUmB+B8ScIPxjgJYDWgykyco96qfWFyDvVb5gRgA5
Uy75xxmjjWZas76cDH3h29BuNPMP5o3ibRuwSgiRrb5AWiB5H1VG4UO2OqHkO7pN
VeK8xszEWi3fLhtr6dmTEPuHCsOVn+likbRsjhTsFI5Lzcw7Zbpz/ZUv8Ycm9+cA
u0SHUZDq9w7OQDa7b1vIRVng4Z+5FgmFow+usUDqB+qCeejWE10IgBgfK0menSnh
6etlu9fEqtsAWHAld2Z+v0xE211A2W5sQxuzUI1tTvxGl58a0Lo4iYG1NXG2udFU
L/R4zLcCh+viR48axR3TjW6N7sUCrOOkvADtbmKpmwLwUDqZ5aQybNc69hcc7eJ2
kSYkmETQrvPD1c7GtQFQWeIxTuNAZaoywyeADqTcqGvyezAdoqOQDTfeOnsIQlJr
eRspLdw9xM4O8oakCg3CzbZ8yrIkzr5WIGQiyf57sXKKoxqz2NXvveMcvlsQ/W4A
wgTxvx36l9AYLvBiBsI0aCbAtXvb5waP6R8GtA7tciU+gUFxqLOJvi6VG2XBhVl2
EveoHaN0zyqWIJRpCBMZ8UzztkPXwb1CJpgKDKQa3XvaZ0P3oK7KCoiJ9yKsuxJ4
JBt83K2sIkSWvADtp3TFIt6iT4q35YaPd9hFEc9J/5HFXE/VwMzspgzsdOAmX3/M
5jUzGO1tROBjPHFacE1kao6KA2Qfb2SRsayLig1N/2m07YAbM+RNXTexKxGcubFN
xbZOG3ccZsL9qVPBlNUFXqV/ID0XejMSTUWdNomwQ/9Ubi1dYH56MzZYNLN7tu9B
RVxWaweNuBOKTmVi4axcp829+oyYReZsmU8Qaj1ThFqiZ6zkMnajUX2B82HnF2wO
3D/Cq1pi6P3tE3yqwxhTH4CdMjdYh3L33ImFbhTH1cYR3mWoKwvHct/MkG4mqIXr
nDaIsuZdfxAPnONmIhFnJ6LVshM8g6KGfWVj0pGdr2TeDCnXfsOLkCjfZFo9whdP
6MpcswtoUh25jTR5efJv5nY4JluTQwPFnh69/Pl2HuSOGXKwdTlKoKJeA2bpEe4h
Hh3DhZpo7gw10mpCBjmtFoACxpdN9CN5UU72bPy6Xpj16C4lleD4jQ5WuVXWHw5Y
uxhn25nqnvhej6TbblF7oNMuX98wuwT+x665RFdi/oBPS1jOekVkwaRbSrD/Gxrh
uvAaJXvTqQhloyOFJ30i+HI04sp3one5fi42XJ/e/Y07SGGzHD3Izo6Ti1GNF/N7
FZjAJ+HKu1PQslOC0Y5QSpJR1ptI7BhHxaE3Bwc1vzRccLcrMVJUNDd7zIhsoVZ6
3iEBseO0tzmN2oMyIEtAXjvu1S0n6mZWvdKVArjdrJNVbNustxMVeWP6i9Pksjrj
Ujp1YKDLRU0Cki0AvWc7/FqFwVXbNI9hXCf+NAQVkkXg8SDjdpW4fdDOSIsaxRBk
/aSCPwtghz8yk9hkVKkaS8NvF/7uKp3TAAfPmVuT+O+rbOgWLgshtTN+nlR0KQoQ
sdlDkY6Ltdy11wb6m32oAqHh68ahoKugp1Ykeb+3d4qsDDYY1Yu0I3Tywzgh17Eb
eavUSPzp/LKPktu9BuPP5K6EjraYct1VE1JI2E/TGxHTzpOS+a7m1qZuvz/AMDqQ
VysdI37TmcpXlFeNBq0E17qm/iakRIiqMhDWyz3RcPmptTLkR1vh9rwET+VLPShS
bOFU4WQQVw4PaRJnQ9bdbEv2bqhtsAW0fvPlm/kObUcRaEmS3nUUutBloXggJdt8
rUEUOMBApK3RE/GhCfEMwKfG1L8B5fOuAorloeamTAEZmMGyJu96ITN1/5H9VaUI
LUGK9jM+7Gzc9eUDmK8gUc3/9ji+3DVgwiptC06n5TIvgEh66/Rl/KdYqzeYFTKe
sOIkNnTwUvN150PNjgFpMp7QsCvQwQJMcfr5uPlDc5FxpzmVIWRLTdAoGqyh2dA2
BuE1k51SwbtUYrp5WS6v9Q==
`protect END_PROTECTED
