`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
IOgKqqFwVZkDqp0s8bTJGnTAFulmnKirZqdJfw+JgkBBZ1OZqeIGk9JZ63oGzXjT
N+Zi8HxtkU6QLtyitQqwygzV5efO8Z3m3Os5RkF2pWpHUY59UHjb8b7QObXvkoS+
e0t4skF4fxKaU2E0dcbWVWRnNO8LhlP+oxSzUP1GcUn/+QiVrwCIfV3xypT6VLHP
TB4EpDriIxLHN8dwdttSoXggLrrWhsOou/3PA5S/RseatEzu9BtvnOxx3KGL0Xu9
tuqi4NNqtU4xwyZ3D85zCdSWh7b8ngE7l1ZjaIrN1MCMv49+gpIba9IPo7lCbGxJ
SDtFeInM5B0X3IM0lLuMWoLU30tp+IYTp3HWPrveCpwdVVI0RoDikRLIBU+fojFk
VWl3G5wuZ+znqTkLcHCYg6nQDuupIa0udxi4E/8Nh6sW6VRfg/M/nHzi7smM0xWX
AxJnOMoPjS1aTQnyO3ffhnv+KqvGreBDF1ohhu0P5uWJ+skFXQykUAH7hpvLK2W7
ptlV9JZpe04xcrPiUkNv34+GJyH5AgqFd/udlE9tjnuja60IFO7yuqGLXpbYSE6Y
BqVANuUXThNPyiNzUYc8b36TFr4hUVLDCx8PNk4lcwtfx7HR9sCtttCMsjEPAFkN
L55cR8LWtWvWy+xxTCgSGY5xesrvJ9R+UxVpWUe61dJb2YZLwd5mGIXFu0MbuyUj
NsdPS14IvLoeOBTp7mAs9y4VrgyQGEVi7LyCv18fEMj7g8ITttxViS46a94Tf/ap
Ao2BFOIQ2QXTKmRB5bUwhZyR7KuKw458RfYRaC7BUc8yYl15NQE0OaeOYcaG1CFG
9pZpN/tEXKRAEJQTi7uzX5SGST1+4UF7frLXfDErSs3Be2jb5OCqRNOrt6RnAQ9W
A7dnwQU4dVNBu/1HDqDiTbETKAGULBinYjqAa/tPCazp5VGGMgHvz3AktP0vF0Q1
2TagYSHS6KiFy7His8J6T3f/TPbDXNQTFeizdkNLH9TpwTU99jJF2x1I7ywk6OEt
Wnn/qTU/1++w2YwCFLgvKEI5kg371x5gJuuI54D0j/rBZKMWcqkbpzFSUbrD/Ww6
K2TVJ27gPEQJfAa46KYkF+2MM/fVT984uZ3SVmE8exkxhRf0U+eceDlMPZELfYYd
hYAgyxgc0xd6bJQqBXoZZKXkV2S6CX89zF5N6fy2lORRTqSoa18x3ZB/u79nlo13
OY1SZrc88Vk7TozBi70mBSooPoEdYgFEIE7nzazAaSVoHQJ9c89EwCyRfEPsCAtu
KBW68LTlaceeNfq1Q0cRLb+p1IDVub6+DdzCJcxnojLnbdmdtZkpbb5vBbilx7G6
a1F6hDXF88cWDiX9jk8QbsPDVOHOo6pXXJsQRD7BKtlXlY45DwwGnJixu+iEJcvG
xygcnAXtigeMldTr9RmF8E163JDEzY0MaB8ILoSgFY4PbBv42BSkAjQDi70y4zil
rz/xfZyElst8B6bv/QMR74Q1DELmyHDBGQsuSH19yRzBBhpcJhE1mbqp1mCExFy9
3us7NR/pwm1ES7N0wIH+xUbqAvYtXDztrIPmerGuZH+eWM8qXy6WPmemcutOKxsl
ZWVDuUWTEynaFNewSyXJh8E8SLVTm/yZZXy7SFCS5Vzc4FdWzu4KP90o980yBBSV
bZOx/kKLPxQTjhi6rHgRJ7bKtmy9uFWFlot/CtfbflgbriDDhPRvDGDwGPFWElCR
OA4mpUtXYnTfG0f+4dSbngOpVcwCiDEr/m25vGApUmv2qElX1JcArPL0IZARJoDf
+LvY56SgkIs/Sx5KpG+MsF/53lhLkiKJjHXDF8t+YPJ79HW6Q6PlJrT7qXVFrjU/
RcQnu9/PNcwFpnXoN4yZuQmoW7IMev6tIr3bYXo0Fd6cONrYsCNFSb4+cI0kUaBo
EQ0b7hPyJH4p20jKCJTcZOAV2FtGP2oR4qUW2ilq06lgWX1hMKFmM0qui26vGD7R
NVjGPQGNJliA5Tr7I/LAjuWHn6dR8Akv4U9Q3rQl3LoMGdv4S0pLQQjFpohZRig6
hKgo63KGBLu3boc4xfx3aDQIPgi+vQHLSdS2UpguTqma05y1hm7ORst0iLYxosZS
aQE6SaPBsiRrBpBC9INwVU+ly5uHFU9JavVSUICCLrX9hCJlP9E0cDRXds8JXeXq
HX02nPF4SVL32J+qJOvstCy7UoU8JZTsbTBvlaF3/nfyM9wnyhtk2BxD1UlGPVg+
/Lrp/K5FGr/kUTYS1bqdRh2vGZT8Sj6xtievQhefYBgA2EPcAf9f8xOAtAxCGICs
Bh1d91u0A29aF6T77auspwOf7J3V0vMShQ0UbP3kKc9OX97Zj6x/8bKXwJ30iujh
d+976400ilQ9sDwCpGAItnKlH52OPNph8iR4uqvZeF7oqUEfFHYIGZuEjSvXE9NO
tGWow9r+cWiC+vR+1HWOTwmf0ioDucfkJ2vpvgSn4bJ2EffJ9OzoeFdXd9sN0+q5
HL+dcbLVHdi5rKntJMuKj6/QJI97ZbpyqaImEMs2KzEFMnYIz2cmKN1iw3jKpWgL
qbqO83GcziF99c5K1nyw7ydXDkMtHkrvIcH6MHif+5DQhukgpMr4WN4dkFrSjLId
Y49yFQ3cAsDGok99PLSoDuTJNUjo0wJuDhP7YS5P4ZKTvjCVS6E4yixhQWXFzNBb
57jDWCI4HAF+cGweouHd2pCogwoFiOfi5tqX8eWZctnI/GrCz8hyamOV9knCwY5L
GVZz1ZrADYZgl2wnDezSUmFZPyqzO1XF+UJAFpSXt/9xEw1Ean4VSmE/jiRkwtpy
gycOuWvFsLXGDg1VX1LWookGugxgtTSYI4A8Asalzi3stXLIn4BFtuYaHzMKxfe3
dE+ahOq7rBBEb1dLZk/gCEQ3uQ//7GHBH1nWhUq2zLkidcBiuGAoMhS6/c7w/U56
SPvpNewb8KDbY6XhhkWQuBiXw8tP5tj5Qp22is4F/FUFKqysFlu4rl3Lojayr2de
C2C/TjznI4zJj7u0AlJVbH16wIPZFcPn8rkBa9bCWzOqhyOTfPwEb3QYc1ttmB/P
A9KWAcoN2/ddaOZqM4BucpcGKGNjzC4Ro2QTF2/ZIjKrZDBMlQ6d/R1BIwiyxZV7
TB0OD+6ysclazkc6GcQe/4N3EieR828NRr4S5l44j6iyX4Ghp7qquqKqO+rc1/XE
EMWFIG9YKAehrIPebWfDa7wOYixTjeQWDC25c4dkWzYhCytzVYUX1HDltNtmSc5y
Eq7Zc4E/HkXoz4ED4e3juruxttRu13ZEenRuDaHKP/B9wYOcjfEJAwj7xJwvxYgc
mR2+soRtgHbdhHSzX+thbPVpIFDVq1KczSEVOyJP8drVMaRxi/6Y96bTvsy6P6Cm
x+KHuZgC9fKw2F69Z1Qq4LzrbnLs7Bf/zSSUaqb7bXpzn7JDqS/KVC6qbxMAdSsL
X7YdV9YCVLFqZkIZwiubL5f2cKL8k6eiOiY1VILrfv/3XjSQL+JNTrG6xnQ5H0Gh
Kw2WlSL+jNOt6dbY/4H0VjIEXpe2PxUXDxyG3pL9KCckOUTAjcsCw4ceAfS3HD90
fE6w5/2WOVhvu228O8ioTCoK1paherIp92p2sUWBLSAGrbgaq+ZniBIHKKnK4IM7
vZJveupWXjvyxle2oPG9ddyC9Hmx/co/argpWh7p1a1v+Nsh1sPKCw43u/ymi+/A
gs1wOq76QiBsR2If6tPacIVzr4SRJ7frIKQgy0JORWW/XqEvMnIL2QRksJY60X+2
Dy7PGpsBlFMKeKcSioQSOHbqJ+HChoeRhYMLkZqLlleBp0HK6oFOs1Yejaz5Nu+a
BUnw2owx69knbM/P/JloWoqoFnf/zmZ0n0zH1s4PckLZFVM+hSxJvn3jgDGreWNj
X+XTS6T60QeShhFqgU6yu8XmcQOinypCqMuhupKsQLxEsyvM6HIwzjGLXW84h7BS
cSxjscxE9dy2ARYP2UpiYMyX+D/gChID9MgrB2Zvlkbyz3BnHDKBHLug95ktowC3
fz5jnswlLcmHqgdFuRUTrk1LEu8rBpAofzScKGJYbksFwfLAe9xxka+7A3rRmuCr
EQW1LR/6HPq/7QasZ33u4OkZ8ZD0hcrl1wXeLaSvUF479ipF4t7inoxrP5g+iC12
tOH1qNpteGjm+yWdCyUmMKR+ucpvUZUsqVsS8Es9Ze1nP9p7SmfwN5mSjDtE7xdB
HZXZmmVTtT7unUeG0zLGVlOIOgsMq9Mh7e5+KAe3YYwaMvdpycldkUoQ5/r7mlBe
xvJ+W+lxJiHrzhJopSog+TNIpcR3Wgo52voqfDJ+IfByvM68i/4lEhC+YsIm2VZb
1Eg5znetyOJo1VSOWL8MiNfg+qBf0fPBZvNdrB4gTiVACPCc8H0Jcx6vcmfu+GOq
Sikzm4lv6Uqac5viGKu1D3mAI8wPAgymOyBlJ28HdK4bwlhOF7uMwOnDDCEJTl8l
TVKFHAsKt7VC2YmriCiLz22bDgBy0MKklESzTpYS1cppjNJZH5eM0WxazLAqCyWY
nL5hNmBY/2Q8q1I1b3I3pGPdzwsMYcmqL/65MqodDNKoO0p0Bo19Es3xOl6tdqNy
uXnAU3lZFHpXAk6asmRR3A0Yrj+j0W3lShg8c5EzrD/AGnjIXgoU6Ee17aMQ8SNc
4uQo861i/EsjFup+9Za75p5cxe7y2FXNhbXrqRmuq0ud0hvnN9B9xxbqKbdpnvMn
+Up5MUSILZJTrpRuT/q78rLU1nGcewmRDWUZDSYAeIRIodq8xECg2suygGBEPFUb
eKsLRVvcFsUlLhUk8lDelo2BMViTFl5zcpXY0l4uP8sy5IH4ixi43pPIlUfX/bZq
raSwVBZ16+LyveTh0X7kUdJg78pDyGWWPF+E127DBz1hS2VgBI/pvdDoUzVDcI1R
QTQs2PxX+C4SgfAXi5b6fBMdwejSqYm4Z/rl+XizFh2JEVSuI9BuIpaz15Okmmhr
fdN3h2I/W94rMvoUCj0kvkLmVhcx8ioF/BuXYYsMtJ62i5wIOkKu8CwbBTvi8x+9
Aje5Lbcb+TXyocsq2V82xrZCc0UJBvgMev7JIzRv259AdR4z9VdtzYe+OvRS6Vg+
RXz52XCtI7YDnBpTL0SEq6jVBQH1BDl+1SJ12T4cQtt0bnbMXUwmMpXxBD17bXWC
LcmAivwSvyRBiumE4zMLnVzNkLAsH/Ljrtbkkxj1p4oUarWGX9xQ6zvuOiUSjssQ
ZMLup261kpa1MeynWGnp4SoxZMZIXMlDXI6w3cczcHX3GVPhe5mzg+Ikq6tVNfG/
3aXCYtkmWUco7IWTSC3dIdvOzN500KBobLhxcUGLkEb+A09SfK7q5znhXnj+N1zz
8Tf3bPJAZcay+aUBa8IzPf6E2cp3BowtGctd9CmpWtzLaTrgqvK8h0Qf1NsVKR1E
u1hLHWlz6FhpTHAbC0PPqPTKOx1z6emu0t3YX3VV1Pxnf2qgJt8q58v1u6P9148U
H8NK/v7aHx5BJRzDoah067gx3Qem9NgBTwY5gvABQR/jBXjfKi1aVYfFnF1xOXtC
3XuoA/3AXyVMA5kwYhFiDUXLHVALtWy97mN4h2Uw2PnOTPlPDCkAMofCSqRLp8+W
x82zIXyUeeV2NMhpEigKKZLCGzk4wRoI2j0jmS30xVjyZGUNo9liD9HsSNkaqM3a
TP0B9wDwVsPh/9bDtAiCzkTv639Hlx4swSVSay17hHOJGwOKvSL8HZ40smVEv9lO
8bNARsNAvrXwaWUSwP+xe4ax1SiVVcMQr9NPdZSyN18ckHxeeHFz7JZe0nMLBggR
JAuz3ANNmXXtxshsHmwsZ+Y70+VfVDnKak/CRqrQB5k2I8mM0vbZaImtFnH58QoV
mAFeSz7Fh0O2W2IJ//hNqy4kEEt8LEcNOo6gsZXqYU9Gd/HY7QydpltiQqULpV9x
T5TWq1avUOnNb5iFTqdyqdJLzJ4a7CcNUzmeRKZYwUVl+0nHNlqO5+h037XCuLo2
VTfhd1Ld2mDJMs+Z9F7MAoCtPxIqzMbydQsDjWCR6fU15fAjmQYDvND9aLwRzqpF
sipwrp19tYRjYpui4w1wIcnkK7P234eBT41WCs7yhhchrerLJ1b2Lw9QOQqKvYCo
ixh21hMEdurJCVU6zKBqSaV4HSbKWqwsRNRJBV1TayeTIk0QSQn7+IcwT0KHEeJZ
6+F4tryixJ4Vp6SDz+pbSUON226Rk7GNVT73D2joOZnpmw9a3kpJKBB4SDinmsJ7
QScL3jGKRftxmCbS6U5NrKAAVFSf6J1JipJnxNTS24wxGLF+f/MthAAWI1vnUExx
KQclLDYmDCA5q8yfibsjoLM3LBFggxzsO/5pLF45rYhoBBq4LYE/xeVHLzF7h9J4
iCXVWQx/tbT0qxoBGq3w+vxwpK6uz8NUDPn6UKsd1oTqGFRWa/gzq6OcFJojDcjP
gnaIi0Xi7Nmqqj025R+SSWHoVXlIDlAG3je1fQn6lOiZ+A628BfAv+HrLKI0Ll+A
4MXlbTsXB9plwKZ985aIc5vd7oIQUHP5zJaRPtyQB8FJo7qZGRuhLhgBPc3xOFzj
PGL6Eh4KV3TvmMbfjT3LBaJhvkjL7xzdulPOpF+6e8Oft/ZECIiHR+8g4dt3/g1b
mJVu6CndLy/SAeTAxg56uRbp+okg0lbvq17mGPKiNjVXYbFVQTfuu2TJNsUzluqH
v4ugFe90cjitfdzYjx0yTgS7V38cgg18oHSlydtdHzrk3CPVjmkimbV0SgeOLle4
pjgMtQNL9RuagPVj/4ahWf/d37p9t7myiOIF0Tvmyz7TEmhx8M7asHej+RwNJcJV
qXo6qmdx1CPfw7YcnMLvVCqzF0ayk3T8Y51TdAcd5BZ2P1+FBjfdBs3f+rAlQJmM
n6tBMBvwhAbEyaDxvHUMjyihp6XWEz8Xv8PQ/x376x0Ct/+2CkbKdO233oqZj9IX
e2BWOV9b3SLsxwOwpdeFREv+mXCa5uzaqhvKIRdmOcgagBwjt7UWQ+jaAfPO9vgQ
6E8kpdtBhaZQsAicCGygQWwXjp7cvqvXk7rO0DGbzvMNL3EWDW8Vib0S6pMDrkEa
250G45HZAPwo2NL5XLTShQUelgAHXKZsvfpNRS3iKLQx2K4XkjR77X5SRq8dYKAi
/aO4WoNAoa/VwLiGKjCto8/m7BmX/AY495YjToYSPDTu640+d2T0C5QHJedLmcUf
2rZcJ7hj7r5Q0ZKtT2fRM+ZEWNTc85LyCCqYjg6RLGq9peC96l90LbgbLLqkkB4Z
SIxBxOwjO4ws/2IhjuhVI8e9OB2JghIpM+691X/3cMih4Tj60Vprgsat0q6ntV/6
XzdvXSenydEJkCwsHwcbna6jJdznMCyLvCC6wmfx/SFnZXA1TjgMcWJhsLBbmgeT
jDQx2HGQ4NPpsj4HDKowGfpbRKnQkjSheqskQHOQ/dgSt+CFq8W1bQ9FVAzHt62L
Gh5dSDNifHGXe0N3Nb/nBLChCHAEniVvzLuE6lPi/wGxzo+0IqmjTTsZf6+ldN1g
2C+nw/riCllJjKwEXjGCsKsk7+zZUp5LaiF7LNYthUvNjwIC3CXGIIGGSOCiQHUa
rEkBdcwproDaozeU6RkaxkrrleiTsqgYzdkEC4TR6Xhd+XbgGQGlDTScMKpw7egL
t7F830F9uWlGGdA5D4Uv021LzmkPTAQtqiEXl08w329rSv8703FhSvl7l8PP6fjp
vwjV9acI6Vr9McrED3bembgeCKCC2eXIvKxxEPbWDg3D3/KtAZ5aKwm/51LiB5T3
gfm0wRHJ+WQ8eHmB/AQwjvJFz1elk43CxJgUeA4iXaEBuJTAs8x5hQBQ50m6ap6G
/0ZN/kWgOpoV+PVLLA30dgRWAc85Hb0hqcYPTvI6Es9Eoo0QAVJRFe7ZojzZrx3s
lAFox2K1Yo8YLUfDye5mdby2FHbVGAJ/J+wRTmoRHBynE//xZ/p/MZoz81eI3kzV
SKCGR9Mxpjj1Xsz2p8MH+a0/hmyd1Y1LQW17lwOSx9H0c0zbN4OxF/cs2qKhsCXl
L9LPVk8ILDfZS5Yp6BxKDGETvhU5ITwr+bLGLrsjWJwNAOwAvsqZswob7TzMqlId
n1KJQni4hP+d3k+AqpIICIc8OApEfga/Kz9f5sSF7n4K+T+hZr91Kye0b5mnYQpr
eomcBl4vumhOKP+Eq9zfVOtfT/9HosYGIfWxSoZCU88imHBW+OH/3g7FinMuyPvc
9nQZxmuA0JbA9Pmmi9OLiOaKL7UTJRQd4Ujd1nTvC0odU+dTkm1bFei8zz/Hw1d3
carTI7Dbe8+Oo64OneunEzWCT0+9I9ojjwiZZazpLUS8b7dr/sujTVfsqbnNE21I
nwWYtK/6pFrwC4tLI69N1mnf2bMH4z2su0cl26sC+NCh6BebKZ4F9UAdmJX74ofR
0XJxqQnS2sCJhxnfRmGhe8tQOsEiDjZ8oQTo9oQnlxP9inbGPjAw/W70Jf8duZxa
IE1T/AgFnXLszi5HhISJpGvpRASCeiCIuoydzEQROInp1bb5WNfRQlRl8wE98sJM
yZ1j1fSQOoLqhWftsYEmXXnLWD9V0cG6fJiG6nCDB6NwA6+FWSOvWyhxZbGVjJGy
LQtFJkT7/y0uuzfQsmgn1IqVG5GMe76tHOq5cLeUjQp866vuiXdpmU1YvrReQpEf
cyWH13WkfK0g60QextNZKU7WK5N3GkFEBi6sUiIwr+P5NR0v8lBVdnSl2v6P2432
9k5HM6dUPao8Ykd6dnzDCaEGZVcdrIOpX9y98W+7t+Q1fk8iICKPTfCmS6nbeGlX
s3a3k3NgEmjxE50xdm5xqyxl3nBSwE4DJ4M2J3BB0bm9l0Rd7wRec5HdhxIdkcPN
dMn1kXyEm17jjaJW6tOk740LfSIoKIpdz97ugyjfb5E=
`protect END_PROTECTED
