`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
NthUEXlwAeaTqAD0n4CMfX7KaNFkW/uCOrJEUS6TSRC1haz5rIs0avy+rMHjlIQD
pMm4js9dX5A1iEo2A2bacTA8NK3k0ji9MJm/zNQsmtILbXjOERpqeznyylatpGfj
Tj0TxiMD5zTUdMHsAt3UJ204zImlxuZ0ma8hKx1TeXyvhxX0fjVNwl7j1PYtE/M5
JkYX5y2YGJFgz7WWQfAR1xnKepOnAG46P8fz5zZUSqVV2fzTk4klyAULmHGYhDPK
z5jsUnZnCBV2G2VUlTH8LrgeKxQuyOUfd03C4RdINj7D+ccM3X298IjVMeQ9syP4
3ZQUSluYZL78VsApYJ0dYtWRFx9X7Ubk3wdAUDomrwz1Sjt4iF8agdRaHuH3f5ZD
oRY63C7TYVvaeOij3r2JXvqZc7j5YLjDXm2lWjW33Gno8Sr2bfwHMA53TZEH6z8J
1iZsm2Bl/ZfbNoT6YatTPerfH3bdoGOmBQUruIVvGMtA2YRorLn1Jl/rwnHQkn2s
uQdBagGZW7TVsJ0brm4ThjQ9CX6Gr6OSh30x5OE1XqfXv9ksLAZB1vcF+WUJmXRZ
qzCNBueAgEt3yKLrLQTjJAJGsM/7Odgi3rFSshuXGcX88CFwX9mWB1M0ONbL+CIL
eicQMhbDtOXcgeTH7glg61Zoo5gL2YjsAfh5gAMSx2FdhH9YN3iVpD1yjDc6ygxx
aJFQLAManOVwpnkI/V1yaZ24vcpwsBSfw/mj4cxTdYcJwO3ujWh1xHywY/vkg+H2
kr1/+11HgslUByghldvAyNk6dWMaW/9zjFU4VHRNOKm3pXDdLWv9f3dKlIdzjVxo
EnoCEOq+0NTeiM6p2jNpTVFPqxEkliQPGGK1iJ9ZNbij0lwz5C8cA6B1lhg7vVxr
4mo9aMlBM697/U5S6wuIzq20gNvXAqZdWIFCMSXkEct9jrxdX0bJoWpJooTAgk2W
LauU86ytu0sj75dwV5lQZzfbEreL3YSdS5KCyhPNU+2Aawx1ggh5ctsSPNjJiiFv
ZvJs383UDeOwzJYBS7X5bIQsHgwmXqYuPHF62BLCQzOvWLd6+sH8CUkWmHSes1hF
rB2aK1M2mpWTlWDICgDYOVoyKagNAZj7UMt1/SsAmpktSb2zEKWitfY9aF850Ivj
ImeMPPNDkJqv9yxZ1z+oWiTvEdxTJsClqsgCsS7tnY4mq2eIiLKVr5Zd4PRDgdIN
rmH0f7SF+h+0aKUrkka7PiAAySFdOz5EyGzsDl+BYj6yI02oW4oHjs7SJgsBjAdb
VNX6WeIDQkUZ6ZmO3d3VgGfpNmhUw6IISXC6nazS1l0apwPsQj0t3gIbtZpBVih4
IAHqTNi0ei+vBoCxc+XC7hz1UWgFA3Ua55p3t4CvwUMlfs6B2yJxFZg7SQ7Rfai/
dgK4shtkJRZncogvaP9WyFgpmfopMBUJPpN+Kl+GmvZRH0vdHQE2Q81XnUA+/3B1
ShSuAycg1dZLQUOVpGTpOARRlhdcq9lFvLgBite91Q/QfpfVbqFMS4BG2DFBqGlx
Yf3xc6zynbFX3yS9DqpNCrBrcTmz6zrpL+C5NQaMtJX7o0HEU78IguqZ6kSJKn9o
lW65cDMYZcl5TThKtlTD1h33EIFLH56S0/iKSpdSPa87Slqs0m8r29gbg2/YUCPC
nr936IvprJuC9URe+knBlFcY4D23C/jf4l2YyP64mZVN80kNhYO6SFqRLqhNWlH7
jbjVyqdzEMCsYTJN73m3wQjGjPHnBEmw3b6K/1KNpr2UlIijzJ0U6F5hFsrQ+XIz
9BR2c3SR0BAyDbERYDC4X503HGlL8mePKAeXMpnnv3FtuOKYmaMSWGVmxkUdK1+E
nlKXZjHPYWxuhhNzRXAKRcVS9fPgL5ueJWdo4y2o2VbSgSp3iuFOOaFPVrjRDqwD
BOOlDdlZ7LAKP6TRSlRrjXmzXSd8mgDaJci69a4rhuxGDaSE8S0odL5ZLnsEuEjo
hsNJI771GtJYNBwaPLliWn+IXuF3B6M+Nh97ToW/SWMgG/5AOlGlYNmt1FXaloLp
L8kGf7Tf4hlXXcMh/ude/4dQaBPEiv65lqvtk0oOsWmeAG6p+rlCDkGCDyqdBivv
ay2Gna0TXc7v9Sp6DbKjK8wqC29tr4Xnz2mmK3Ao84KbdAHNekBqOjVCoYFz0kIs
ThLYXhG+TrrZ0HhPy/d/qo04c1XhOFPqXu27WiJTY3Dsj008gX0u4BV5AIEf/S12
v646zyvxwYCVPaOYMkqkZCJcoX4ZfRfS/heYJWse31N8ve/gDgtnZ3oy0JnTjris
37ifILkYfPyw9FTObHLrUhEHsP8SF50CT4Fiw+D727UrXXGEafYcFJc8v0/Mq1oe
xE4Ni7SF747hS5XRzab7UMJZail+2A+H8lRpWVXojNdCdr0mjj+u7idEXNLN/X4+
s9T7on9QCv86lDAaX2CzAaS+MwZpQxpWOBVwNwiSyLdnD8pl8zDlto4l8Qg0qFAB
pquV9ZC/dXkE8xSqm6RfMS+3b23hcxT1QZZ0rupcHejrt4s0oL4MNr/8ejG5HyD4
P96o9hO+0iCaDT14V6N1wDUySKCvMOlGRdBN+OaUJP3kJ3wRjCDQnglQsf8aMU+X
4lVEC80prhsbJC6ejNLNzhGptPLpSfSPsHx5xDu/HB71Dat91LA0b63bZWxvepZ9
XZ9XO+AXvbPvTZDZlRew3EYUabac+8lOvD4Tmik2yMhzKTjXjZME4tP3C6Oj2vFr
wwmzyqAvRAm289IfUQphwhLKeugpRuXl7tYngmmcfZXtVS5PAt1yA5P9vVQf33jF
cwFZrBSyEqM/6wM8QfaD+xHXs+rO4hu+xv2s6KEMy2EKcauVYU1kMKm30gU9eaIV
hj3dGLAIU0/vLN0xk5f/Wr/mNluE52KTvMI/nxWxqY+lsvSx0udkXIsYamoCUFsI
MY8cE5sYlo2B1on1KaPrfXLiekIGcRA1+NhRwH3MisdVAJ8eNCMvZwaLVZRlMGt4
0iOSJGCcYlFuWaM34CJNBswywctJBEHiR9riExVnTrl/CZSrXKU2dbPw/GxkYUwO
WHXZMTOCCOa0dvyYvT3bpDk55d+p2BcxQqpkqnP/Ywers5KWkoS7vvkBBvsGrd7f
bZepGiS2eMQSFnz5I2jCUItKkdgDW8mddg4l25T34oHhtxuyPjKZjgz3GLTq5RXz
ZFFGs6lLkgqnvRXNJBjba5FvdRcilLbzJecOl1ey3BgOejaVhUV59aZfBItw8p5v
PspqNCoBNcJ/2siZ3IgcEfRtSXrij98juY53Azc1KeUCzi7p+uzuepHBDEvKLST0
CTIFwruO11mWh3u/wdIMKTjEcERYKuhj2B6ObgIKiRNi5Rzi7Plj6sExEoLeAUf2
X6tFcbp+hgr138+sP1K3X3QSm+ev+Ibj/h/UdIVgJChMo5ionkFAcMk2ipFnMX7Z
ozGESm4xFrX+dS2VXc77Fs9ttYyaKV/BIHf8nRHRqaFeOUgTuIrglhyZ5poQbulO
MS/aCWhxhaG5zFCblunsbFpJwIpgetjVC1+FM1qux2dzKYWpDI1QHdFYbXWhwnir
Ip/092hWRf7Ai2bPw1Zy5wc/vt60W74tlkCpeJNncHkjQ6VZWnFgqjRr4brNQm1z
bBelQOismb5VEjPr60/dIeR4HP197HW5zSsPGwnMxrSQWxE2qVHX+sctSnLqjYPJ
fv+4nV59S1BELOsOpVgrAEZ/K8sg9qspCZFV6JJAfX7DHfuObNpZAtR2epfzzhaw
MVj92BviPG2/7/hXm+N9fpZcxfno37SXOSP3D4AEVSFpH5/IYPsuxUUn21TiZkwi
j8SqHPrsqvJxqLlrLytYLZ2jyzUdYrnUZKttDCEf5JbiqBhfr0Dy9FZ/eiuijpU8
0kpU25bDZXe7D/RBYZ7SOnfoUCmjlE/kGKZ5qswuP0dH3NiyFv6TCPmGHYHYWNA0
dxiDJtACz/dxbOYInHcosqh19AYUf615KGwPJ2AskGEdYnt1cpL2OfrCc3i698pj
4Zb7CLEq4LKJzZMFX1bj071S16TLoUKZkRbtqM+q0OddDJpHP/SOHLWtMDK5v2Y6
qXYCV+WG+2pK2TvPWw06FfgGXPOZhci0pZSaerQa9lEEXS3QbzkyV114oxuFDyJp
aSzqe64OTJy0UWAbvcsQM9axYdYX/6hlFvSsemcY4RVpwVC6qMAAvz2rB0SiN23d
28m76cnjqlDuB222c7TVvwpAXZJLxfCsmH1kR6/1vxMLAKSLCOJmMgjbo18VsZjF
QW7H7ozpOYY0NXiCFvJ3SzX/Sdbj16Brw8P2dQl6WlDa/C1nHQuhUnCYjlspcyuj
fmNxtPvdOGULlh1RV6YuY8xySTslUkqFLnLuILx0rWKHP77IOjf+hsFSlJWIYdR3
BCK4YdqfImEnYc7h5RT1B7w/GJ7hz6nL5n6AcOmAJlnHTcTdcM/Oz3OAwwuRMMzX
i0TEDoP2uNI/a3pFn/81QY0NIFCLDAWzg9HvntwG01UX5czuYk/5JRaAPnL2S7c6
RPueZChGPIGJnXSopNa/fs2EQ/117lMtGTszaPLYcYSEHj8iZfL1htKFSW12kbvW
M1YmcnhgbpcgPm98AtKj/AUqgOfnN0b0RucJDzqE4rwfD524jUPphx78nKO+eEqB
sHgOmMt6x5rSc8YpRad3NmdGkbuUjVhSstl5GKFB3OiPH8w12QdTMM4mUbYZty+m
qbJ/Fmvlc9iDGro8Vk954cxjz7O1Jhxb4LfWBJcXqpPCcnpf4X/mJCgMtWbtxDeH
JxmVyxnDwIWK8zfJwEYJ9m1UeUZ+W4Ep778AHqYeDpr2SsV0yz6uuQnQE3lovy6p
mbc8LiZYj/7rqQbgzPyntBaYSvisZsZAeuyFFvY3/Vm42H3eHn4faRM+ONlAzQlC
E5aypQEAZUTO8xtDDZQ7pNRzv/ndr/gcufO/aEhuHBCqFEC+uhjMxX8YyzRfrN29
0WC/QQxApXsMdPByUpkmyUIOEI31IQz/np4FVAFUIlOCT77GVAPLUK6iuDUR3cNX
jssSjpehiznf+FcZYhnOSkGttItEQDC5sJgU+zdD0erRk5GS8hcMpXTlBUpTEb2M
V7ML7BQJYSbzXpaYZ3+TOZzS7thl17SPtwbIcrc2fGkIiZHWE79zQJSO8hXfFkJd
/rjebcNtwv0CI/iHuyevB/hf8FWwrRMRg/LVS/UnaJcVJJV/ObcZEWbZrkGQBYYc
9OL5A735wYYgeX3AGgMbgBoZ2a7zW3x7PuC+CdYZteUZUDn1VEiut0F+d+Iu9pBP
2MY+YnK2BEWWNgynhPAuR5YG73cSNsU5SDLQ9nSkfPGJQZKfvTCYHoSxeson6Wto
9j5t+MO+phKn1+3taGChYGtKPMuKg9fPI+AyBpdRejt+kJyozFVe+o1FghpCbI3Y
mO1Lv1gl1ryvVJa4pZKU/Mq2M7z2SCSbwRA2qn0JJA9E27VrkZ9hOVyuGs/GwaZD
u0Dleyeks8bjJISk/hKUO9LOs1OZHhP5xHqMqC3CC+26CX2G5/Dvx/ozVhBkHYzN
haPpf/Lk33Viz08KSjo4y1YewGW6HPBbPc/8MQ0ghMFtPzq5IKe1fHBzSpO/W9Bj
B3bvZevDEaMNMz8+bG/PHIMt8UQWCICwK6S2a3ylpQtvg3UGKrSGl9NhU75tzp5i
zrOtjEvWNO5qXMPTJp6XMgBdyGqYrCXcxjsQzq2eHcpM85yHVv9zZ6a2rprbGEJ7
7eXoioJLvQyGwGw/+bUDtX/I++PZZlKeb3b6zdqPpr+BsSz1yeX3ckXx0EJwUgb6
WrkQU+MeLRa4rVqIEibLp+Hocu4XVyda3y5NBMP4O1FNUhtywZGUTSKn8gdn+v9L
sP3e7viu6/8mpliFhkrDy9lbQjpQyCyq8Ej2jCfR/aAM07PYDLCBDaUQne3OiK9u
5b55V7j8H7NbySvDWH2vYnihcqjvwtG+UQEptkMoADug73DN8+dP/8K+fq9lRQVr
y6ZMkEVvyH36z3e1ZpehTkrnPhd6SkoL78bHtenquD3Wy6MoQjAUe3L6mQkAjYno
Vh+bWYugZfFenJc+33UvmtOkNb8bj9SZu+Bqny6Wrfhb2Ki8Jy9VOmFCsU0VcwWh
CSayzh31x/3GO5y1FuVsZuSaF19vQpKPobGSRmUjnDgbZb0aPm3VCFjRNTGwgFCJ
4VfUg52WFXCraY/Wj/ERljPijnSHWtxs/xEB68kYfRd6r4TzMDv0sV+j9IXkAR4H
ViAX5tUa0+xDR7EUKwlMzZhcCxE6LZyKWe53FlCt+RUxQQ2eM627jgmctwBHJzae
dvo4Q8/tmAktdyZBJi/IYazzmigMmZo5XwI6GDB4ok2haJX9URJY/nG7+4nyP6Fc
DgnwxDDXO8b2Azgqi/ZUp9w25IqE2zb35+l1yZqs2ssR8xMnOKV7Zv1S+Yv7ttIE
jbF8DYt5E0nBLxHTgWAtZoQy44qWpzA29K6YlHIijuVdIg9E693sOUCHL2nbmA3P
iqUMzLrczARujykDxuAwHf7rU4Vgo2K8L4umS/DbmowBM81zIGF9bOzivdPEV4Wj
xGy82BwZ1H8t6h+oihrk1D7mIcx45E7pRY2izM6e36r6r/6eauxePhkVuI7vL92Z
rg+ca2+aEe40fycRu0m8q6aYBbz4yyxk8YBN/lvG+5g=
`protect END_PROTECTED
