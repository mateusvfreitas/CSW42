`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0uIll7EjzaHNdtBmQTCUOtRaMgTiMLVhvpRoJExQRjNwt9HYhnW8VqSQyJpFPECt
0NIgiqpvO0pBA/TxLL2ObWUJSBLCJyaTydv3pzcFmtlhlPh7uE3JNZgQIjC6viv6
0p7Hcxp9BTn8I+T2nZ6OsFK8Amx5xdyWgH4de3KCDb4AtbZonYBSBrIE7ejoz02S
tATNAiLWrI5GlL0l196R5u+2dEr28hyNc8rxMGLGJ5LezEkwsm20v+OTsmnAYo6x
72X7G3Q09NV7AVSeZAzGuzR1wBSc0spzHQ7E5+nW2xp8KeAp2u/DaZlcXxHWZtc4
9rH8tqNIakDhdiLtYIkX0FJRfXIwxx77wW04vTgQG9jqHmRvTc3Gj+p7gWGwV/aZ
XHN4IFboDMFugbUFVHsOPhNJTIIkiMEoInEgSUUwYh7QF41KYNEF45yacfwdH9JR
dwJK+ebqzKIF7E+I97PjIDXCuHpuaxDIdroM0WiSsJl6lOHtMP7jICn+TXqaMsPh
k0tB51zAetytJtJk+zO7PjjoWNkYkLmFJjs3QZ0K7/eS0DAm2i8jB/+2mxeq0N6Q
QexgYSpuetqzKl+zZ41ZuS9R4SFiuE4Fbg9yc71J1xoqgHnOwMlTWB+iAdF91Egn
9Y9gJoGGSRLY0s1K1/RxEdg5rp6eLowU0XDifmZuQXAYqSh63gT3YzELDY8W+uRw
y/2v74CIW9JBy44RJckIcbflNyGYiUzXUYeuQKBA9cPqLv54PAhFI2sNApTe+By/
dy7BNvM8NK+YzwNEndUgZWJ+iOFvbeZl311J/SxSU4oVo97GYUGF2/T7G0mGJSC5
M4fxTyEC7ER74TcTYClGKjgiFcYPkbkvyagt7OrufabB8k2wbp28xtGuN/1ZsSHy
g528eWSnzvsLYLmti3B8P4WtzGaKq9MVlnrR0dk4pzh+8dNf4uHSR9gMU5eX5GfJ
nKtVfcWEeYBWRq4kvfbnlP20dPWiwjamdOzixwCKvVoua1hDWOhtXCACNRb/N6zR
8IkdEKHdBnnYyYfiSyFHEldR2nne5N2JD/QGCRpWL3qWF17GdUFzX8Kh2hrCOtmW
YHeMjO13ITQoRrkJ7omq/Nl18cls7Hzv06+pkI9OpV+LjzC200M+3Iysa2xHxLnl
/x3ChopBdg8ZfaZ+v7KXDSjCmO+yjom3nFtcKEdD1Ul2RUJrQV4WTRN1IObQ3T28
ntORWZnqtXabWHvJ06dqVd9tqWaBLgRw8i2/iHnQPq+Ys6qqBaPFMaQio6NXio4x
TDxKXUe98FwsaXWwv6At7gaKdfejIsdGCweUn8gORhUK1uNxlwH0k1PT1UeaKS/m
WZuEMQ8ashZqkAbflQ+M8LN2RI2gBoETC+JH+beBl/FBEmVd3Jtb9b1ch39idpMv
ac0DoDjLOdIl9YkPYds4qVt6AyNbUePjdLLFQ/6rczGTWL3kMdIh8SLIkeibA9Ei
K9SPrv5Q4xWKzaqrD7t+R2cGO7YzmZPe1cSE48XZAwcqlYqCIQB7Us21cPpGwrwd
0ZxPzb6kewAp8W2rp4/DNKAxcF6ITeOz1/ANDKuF2adg2XQ/7vTzAkxzsX1S1kdF
xe1Xi9krgO1X+bDJ5FevQ+HLOq7IbYz8jllp9IWYqeqd6nOCMyQME84dUZGOyWG1
BZiAy13UXMkDb0XV9Yjf+H/zQAg3t6l1yH1dkFOKgNzUug9jDBo/2X8lzPr9Dxfn
ONYUNn9KNUwLlEyiDA3lwkTves6hkwRFrTLOAk6miHp+vUlFYn4ygGLv6GvVKCCq
nR3mmPea4w1ZlwKJ/vuEciRkSG62OOkwv5VKo9oaPH+mRvcQiKg1fCNjIwegsI5L
Jq66lmcATLcbcOsQb3MAZZafPZSRlxVp+H0znFfoBOM6WDAn5RE8GqtKdaTMiaOc
VJ+4tSObRv6mR80/Elv8Reivh1ojm/EB2TiaQAZKTWjlAcRyjE2QFmt5hhTypcPT
C4AtWdp6BW2P9Xrp3ea4HUE7IbKWTqLop1pfNpVaSSM5wyJ+BUywGvWyaxfcOPUa
`protect END_PROTECTED
