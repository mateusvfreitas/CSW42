`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
3hTQyAfVPja6p2La5lPB9UNPlFrg/7j0c/WBgDOcu7PQfErgOq3nsAHOQtyJQSM1
m5mcn6a3aHv5bxfY70tHjRfrxuecbd2Oh/a1vJ5t5mIDK/nAbAVQPsTDXv56YaZx
pq5qXTj496OxCR1XXwGSbbVeUbjZPwOBbLkPHpR1GeFQEDiGA2bwq4qUtgHg/4RV
UhQMI4a44S6t83COLClITius8u53DqMEVhFDAks1qi0gCGAqZV4njASPw2dVwCm/
rprDEOKcOQrahvJMS4RBEt6TtjgstfTpW7OH02aMo6FVXhZB+Ft1hhXigqKhl/51
xv1w5FCEkPeu6ccqbp2iny2ydSG26kRmKLOImPHo89WmCbRaSA1T9O+d0UQP5OV8
SnT6irAXU9AP8s8QCMF9mLLXar5qQWwIpMcTmusp4pkbp0Ke+MYTZzGvDT3NLg+9
U6ckvCZd5dO+KW+WPz4PYQrB3mQzYxxUBFo3pVMqgHCRh3JRMZ/VO/sMY1VxK36o
yB403ORF5nUNfnj9VIV82OI7ViOT+zW3k4lrhxyMi4N/nDsuDsXsOPWfiuPAnOwP
5VNac5FirI3ZaOoaWouoDiZtgbETeZp9pffqFoHzv3s00N09YJtTxF1tnI43E8KN
K0x9IGkby2Om1LrRwfIX9PFe8/9snOwUOYd5wTynP2TRFLOi6d7bAY1nscRV4DAP
KLWnRzKx51EjxiRq5M7QJ+SQkH3ceQlqjKD/p0BlviEE8+UhCywHGijds/Z84Ydo
0dLKh2z3aPnuqiAobbg/xmNiEsoggMJkzEulZoIx3I/oeerWNfQOw/PEEwZOnXGv
A06Do+ZUMzHNm0OgAaTpmqD/4OmsYfF68+3S/SDJ/iVj44BUZzDtx1pnnOh7zRwq
GtD1VWMMd2PbEKryHjua5sxJI/D9IOTiiWmGTbstPmY6ZM7FHhBk7HWcr99q1gtQ
+gyJzwSp2P3XUM0A+onX1b9bEg4ZFMVqJAkuwTuGCNpNZ2M4gaK+Q0lcSUYDKlMy
OXrEU2hVT5Q/yoIuHR4WNtOuqraiWU/bL9XRlmQP91TotBxi65q91OmFwlNWwrZs
p2/xlyCeiBmN0yOKonOHupDhQS88nn7zLNnlMjgSXSIzzJ0S3qjdGj+3efKiVHeC
uUZ4vOQ6n2SS0gWv+IXfdPNhnd4AMJAZbgngCwwN2y1AQD6E/UB9gmgPg75984fG
EHA2AJaGgRDehF5JcUOpRawzuTWec3hgNUDsknmBOHuIVQscFvBd+Nyb42A4yXOI
k8CXIwFP/N64f86YRTv14a1Ur348/paGeLssW6ZoYHff3pKnYsiYYeM70L3lNXp5
Pq1Hrrnz2UCI5Z0ay5SpqMICcvaiinNYadVrqAovSKYy5mqP47ItIAgiTKiPRSuw
nq7CKqKLWTTghLTQKjhTsVTjMhqABb5VdgF6IsK4d/SiPir1QXj2yoEEmkHRlQnL
c0OE+OakkZ3b7HmEQAaKM4RlP+COdkq1dhbTyIrkb81npsJlvlcjDF0GH0ZyWiNV
oGdPuEmnHkT79n3j+25+c4uzfWRiPlYsKQ+UvZO8rKbFvvtOcZL9ycIdAiVl8k1E
907pNTaab9LSgxIlZ0s23h8d5XuUbxsgOT/GXU3iqwrUlf1xe7KWUlc3/k6H9Y2S
1iZMsLmYuwWHN2so3VlWPpGnjKOgzNqOpu06u8L4KN50PKfz6x/W+ecNKIKfLNJx
Yh06I5W8024GAaUg/n/p4zzW3Em68BU16OB9DRdk+7Hiy9dCbygKoGP9wbL8BXOr
xJujxtqikqQa7LyP4qeTluqMZu34NudUyLwbl3J7aFl7hUTB+lR6pejeUtidP5sc
6WABvi2js37lxSwqs6NNo4jd8o2kKzkg+186r9RPjsWcc2DJYXBCCjuyBk78LqgZ
dbs9kgfTgu0qjj3H90shiFv6jeTYH5a7d1woqusvZO1i9vQ7n2WjyAH7AcJeaaDB
Q9qX9qzlL77fxW55wcqKJFH5gubtsZkJBXwpB7F5Oabpe4WQyQcAgyJpjTzeSBl2
u/pnyEI8bIAZ677aF/UNqaZuTv9me7zSrH2b5p1Sug7/3AewrX+Qgopi2CD0YOTV
5p9awp4if1uxfEIjFUMqZjyOq/vbsQ7BUVMwHUeg+OGPNofRzslaRRZxmmp30Xnk
yezrREgxLGhw75fuXKcWbrbboqoEbjSNLCgXZ5NIHHczHR16mm5+Z1SbwSp4uMWR
WVj20KYHp9dNi7e4dnicTA==
`protect END_PROTECTED
