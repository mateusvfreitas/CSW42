`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
q8dzFsl9XcBGGqbUwNndgwXZdpicKIjrmry6zUpa8kcVMRI681dYT3ZHm7Wl1eH/
Jg559Ww+/4dV3fRe0CBIfD6xCHibJxWjCL7qz2uw3O2eJmIwmjek5tgXzA/aDnXX
RVYU3gIURSyL/QCm3blrCNSRZPzpmuvZktY9PAoMeyAUqI5NbpcGRnq1RBzAjjGL
ktyy3lKnHhVPk/1uS5U00PzC9Ao6RS1VAJncD4aPnDDrxTS81sXSa+R2AdcgbeMj
K0HeesCfJF4hVceHe5hEy9AtJCyYGl/ERxwSa7oaBFfwF39mDpUgk1JusEFFfDOV
G3Vu8xwMCCdCvAbGTX/9Q/9DLf1eOB62jJ+m5SY++izh9f7DKAdRqDS+c1NPj2K6
xQ4TvSnvtfe54oJS24iR2DtMmkDvqplszD8eClk/ImUQB3HpUnnP5wRDt5tXEK4l
6IwQOhqkweJce4mta2oEBm94wsu+L5at6/56m5AnIipZFZZdH9htZ7V3pHqvGHhY
yKbN/5XRAn2c7RDcEN4jsdNbW3cIW5SM04CfcPerqwCnl4u3Rn+5Jm5MJ3SfigDz
HHgAMBRFopc8YxcwpT4CFfTcyX+sLVTWPDdXj3Kho/Eex6jP+T874Ma9tOidhgqJ
mX/aHEvQyfIOq8Bu4oOvk5EYmy07LXcjLZJISiuWjqJhs89HaldFGMfw3GdA41oR
hZo730t35c0SswJKkfxxsDaV9KpNBNst2tMpSFOX4ack/BmNSA4arCMH2CTZD+JU
Rn3dRMboRpvwafd0hntHPeu7RCn7a4J+BaiaTvj9dSH288wP8ztqM8C2i2Mp2Dx5
hUAXv9+2fY+NXy3h7ANNPY9Fe2HYw0wke3Y/HEsSqkX/LROiTrYgkmwRnBbxe9eP
Ujc1Wv94a8V1p2EfOKpJtHAJ+Pdm7nw9sl+/jlQKuxkcKovaW+0X4KVNg2KssS/m
4f80UgzvYOAl7pkIxn+vb7b895z+2Jq/KWzrprIWG5+l7HGo79Dza0tY5LUWlTqm
EWmZHiQMS2qObIK3rIZ6z0doN+5RDwovg1/vMWYnWM4wgRTGiFTVfhYSISee7OFR
Pj2uP1SkXJgGQIhGFoXO1lDIsJK3bZ9VkYQFoSCPvWvrybp5LU03uJwL2uzsVAW9
P4WiHgfhytRrxG4yFgSm44oAWGptfwI9s9Fgefl8vCtrxnoxqxS04wggh7dUjf8w
6p7ohSHQ+WgOX9OcI566j0la4xVUP8oR8/WR3T1viIfQ0XVpVWkekwYJdsRW/Wfs
1aFrvaNjTSmgX8HHA2XoQeMo2azBZWvndZw4of+t0jlM4mfCVQyV03hI6VsBjm5X
CLGehNiJ8SMXlBp5DUJY1cQZaS5od/zZ1lMLHHDWGgcbEU+r1IA7AqQk5HL2Unr6
5U2YSmrJs9daIo6q55ZDXE7QBnZcexG8RocGzl/vMc6R8PwLKL1vIXjhSNgGH+64
EOw9qpW7bjEMy8SjZXz8ZDvaXRCWC2hjhWlPbGp26UebDQY10lJfWKNINsjzq5eF
gA/2OkwysLHpw3PjNEHZjmVB09KeEO4PbFqZ6Tu4Oahp+Ct6xY+awPYirsA78SZq
FQTwV004lTJtALxjrclHY9Bt/8oaG0QgbVPwFvkHJZU6zr071tSYZxZNCZXzyMlk
ID+hSSi6MFi8ibJ6Jfnu/zmbBjlKebdtvCu4nvMrBMVgj9G1quKgc0wm0l8+1tBQ
PSrLRrhNZ86PC3Sc34YEPjoc00QzWU081DvClVBRYbFveKGjYHhkG22l60o/BsNP
vW/lSPK1H8dk4u9uRjMEv1SKz+T6RsQxjTWnVy/rTeM8ky75eg7yjm2h7hh+fXEr
qrLhsEQmOFA7ByfJGtt5Wa0ktB5JYoSZi2TLEz2WsxaUI2HZcinjoI/uVwBd7cv6
aDGqPLMYtGqeNoTP6HHda7KAhrDDxzZ9tzOOIK3b1pQNz6fw9nyhdfWS5sDSyTHM
o6gYp7/f/iza24XcAPGIOqHLR/Sa/ioTLLrOnnJuEcvzpGHl4BM47J/PezXSBP/R
D2X7cwcdjfvTFlgIuv5QAQR8O/pqq38Vq6KGxvnHk18aQKyOnbqdKuDnB9LCHfhe
+w+ZE0s0M/sTWFJIIYA8CB++uFabSokrDhPY6a3IUUPWlG1J48oJ5oRjec71Zju+
WC3HHXCGfcLe+b6A6uRKaqyVH+PpaZgbgpX4KuJhPh2+F8tnalq3nK8w00RwqCzu
F27Haf/ueAKuhbq5ihv2XQbv5v90cP++nzzj174ORDRkaq4kiGlveI4a45/j4OrP
KNmObl+hj56VGy/5peSrB2T+uSSKZ2ux3DjcbTRI7Ge4bpQSsmTrkpIpwSHjTQkp
H75jzSYg2rjqiYBNgcvFMIyFaoLTjt50DBgGkx9ySmvUikCWR02f/C94ePPmypJ6
kGSqqzr224g3ZUp30RijOeVTai3chOQW7eFlF4YaYqovWiPruFZX5qmiDV9izUOr
N7ELNekv9t1oASlu/BgoioD7dt0lc7ParpFXVFqV4tOrlE92mxoz88EmjhJm5WRa
AF9wj3N/dGvlVPnRf5/hmsrGf+gksMHQ1F8TsL/XhWmulS/dUjMqQOVu8rJeQhSp
YH5Sx4nz8yQaMh2cFTxxs72KcIrAGowF+gLkzquK91CdooNic7rKKV4Cpgez7nOR
1PCiRP/tIQUnA9s/++rUhTz4SxdAHzueJJ98ThZ6GozAnDdYeSuiC1Y08CXZaL66
kH8TgpCbRj0N0u0T5w9ErzmeHHOc96x+cThqaUhnKq8oysmBKjDscgMsGEL0/DJn
GglddvtnYonOVUNusRP1b08oybVZxDR7Ym+I3H2gH6WUgD1LmFApJEX+8c/av9Qa
thkYUozgrvO8oNpuJwsOrbqhz4J7ODtYzWcT3fNgnY9JIfQqi1EnIxTd9HUWN4Wh
cuuMsw+OXqHqIdG+WJSMQOF8sZ8AL9N69zRyu4Ik5dswJ6mr9LUZaTcXWwQVxpO0
CSu52lTXA5ue+MDwc67MBRgtWEvGaxQSctUxVmfurzfm3UZ5okVsoDoJNv1aodUW
HJ4Q91iRIB1+shKAWcolAq0OFbIbXnHrrjfx0Oa6bNYNxdtHF4pMLl35rt/mhlk4
uXB3I2JAQZvhuIbk6rNJgB0WdpqggOfcl5f9UILh/kb0Bb9j44akLFrbFBm1uhSH
LoFBMFm8Pwa1y6SdHhotag1yY03I6wIpljOd3lcuLvkqzi5qxA19N+pvaStpm78A
Janj2K2h3riGLJrFYUMVPPRor8w0DCoUv6SjOfkIKPzUPseorJ9WNHYyx3WGN1uR
bcc6ccrW0PHrmSPG4oGXUkkD1CjE9snAwBgwomDYHeehV3uMFftVvUMIoGPiCDsR
tfEPzUBPf2CQ8TDSJrSLqBdVg9JGW1aQY3+7nhA75VH61LU7hT4YNnxc21LpaP9h
VptIkNjbBubWax+WbqpPi/SvL4/ZO9zAbm5X79Ec1sjb1KtsLOkVM7C81cM9DIWM
kwZudq8wQ1BN5k/KcAitS4008lofHucQ3ALTUxZ8k+chMdc/ZCFbWqMOpRDyMemK
Icow4iayLI24HxgEsZ6YxPwMNBesiYTdApWVw9JPhULZrtrupjP7YL10EjvCTzP6
dgxT0y4V9y3VE7W3L5TWos7yDGS2rYnNxN8aiWIKmJQPe4TiSPBvQ9TPPOoCBLI3
sPh+4xqAHhkkSbCm91DgmAzpT6G0OAKKFXUYV8+J1vDy9+3mwmXNSVeHESA5BC7O
92Nrq64+u9BocnmvBXote/MdNhhLNggGDN04/AKdpyMdO2NbwExMf1WBU+BRS8XO
8BfGk4q2OjIFuREDK14g8nSb100aDP+aE+fTNZmAYP817qIHH9eNcuCqe28HhMlv
Ww+ZCiYmqKPLnECq0vOqedGHQOQT9FRblpMfaQqscvuEc/TkvLkIaP7r8QdfAsun
MyO2IP0eXRlDi5+HICc79+U0V+99FgimYtE/saAKMM6oC4du1W7krQvHF1LxS9HD
+wmJpp4klpdbRNistSPPOgP9zx6WAgiPgwxzpqsH4LsR0bdapYenZnNIywxUwYh6
j6hpI4TrNgusilROy6MlDFWdK35AqNtWeLtiNj/kF5JQhqowQ18LXegyN3ZR95q7
ECuCOcZ4u1g7+5QKMrLQ4PgqsvDD4efylei2Rw7Y7lOyYHMyk8yMfC43Fw60r5ug
a9TJ/DaThknFo8eWFNY/h4r1t3r8gQuBuVKiF0N/LQ07U539Tad1+l42eW8kmp5A
e5rVTFoRarRWkSsvTI1P7OjzNKSsLeH7Z3seOAWOqxIj7/zRw3mb3ZFRTtiwGvQo
EALNabQ6yd1zcksNKaryrD6WCTPKQTrGLJJ/CxdSnOhMFMZf5lUgLtiuLxsXwuoj
fXH6x7TsrIdHeIiIAlRKwIFQp/2iI8vxkJE28WxBL1aXHW369sF1vrG+Nqhiq+dh
FNHQpX4XmnV5mcULgkHgpqXmgj38GAeVtdptApFHDhDOVxdUxIY0eiz7/LayD3ui
d0dr8+OsRDt1X3B/vnmFF/8t3SuY9i7LPRNtYHXaUv/OaqmRXuHrTkxjil8MPSV3
5huRZzEcVxA3SHo6CueqzJOcbsekZJS2PbCX7Xh2iY4vOdQ0+iuO0hqykd4gYVpW
0nYgf1596T2dVIXWAtYP6U655YYONyxDjWZpFWer7p0cVfimQt3sCaGwHgJlKpFH
94J4dyK85bEerQzh/e9YQFPcMtRgqUbvKMtNmScm2w5HzVW3YB65aO1Ri4su1cVN
kBm9L6XvorfRSrx9KlYwxdBMzBqw613encVIUinctP8mN2pWGJLG6u8U6zyInO6t
7a55a85tsseOk7Xm02LZcxEi70fSyReQ8iuL+/R9jHmILFuMmyatpkq7RQFPHVwl
zBsiwnJeI9QqJ7kAPK1LuwDj+SmAXQgopbyyLnaQBhHpXp8AYGSQ0WXhhUjNZOeh
4LOahKMLcb5OE85u7wFbX1IhqgXgxlsYQ9CAExjmxwqATAMVXE9M68Db3wmceNcK
AhdELAEuy0PSRXzYtkHJ68A1EEqE9h0k6XBafynADS4J4rnHxsHsf6uGNNsfnZfP
sweXJrNsLOc3pjG4j1C6uq6YNlVSU786RvDxxbUoKsyXgjfaR680K7dCcI/hH71I
bbjL/3OOuxk42ymXZ+c0UK9twmtRRiv0flTP0T3oyJ4FkgZ0ZiTk7InV2+B0Tlmx
UljHdbdJ/S9NuOHmh2jy6nlivPb6CCk357BOcpx0E3upBTGanes7AJttM2I4Jhi2
ijoPDtz1Zjtd+tSroqrA6B8EhcxBnbG2p3bCCh9xf8MTxJLHCstasfjlpterEHXq
57a7HXAuwzDzjX2V5yJBZxSAVyaAPOcbnf8QCbwj4HwVhkvf2KA2OSqUcOYgd9jg
ivHowUyb0POwqWl8Ct8Q9c1TzHUn2gSv+EACY7h3XMlGlQuQNhhs3M5qaLQoXZgf
gr5UFHsm2207tOkWqOUsrR7NhgMZM9+djLtuVzs5BvgFvGdPNZJGv4eeg29qAbtr
VgVwbEB2wqSWpgYGfbBmF2skbY/V+ktq98WPD4Nc1TEUi5S5FjvyQ0wLN/KxU3Ks
pPfQ1IZ+lXOAiBkaZBDwArDX5m7Z4nBzzNLDvzv70ZcF1FxeCAFrjcTtbfJCkARD
Bphcz8wu5LANDLp5o4LpYBBLzOPjQxFRfXMc2EmHrtAnhUKiN6Nvbrq1huYVUiW5
qvE7Q/GNhc/WEWMnCY/T4OCaOqap4iXCV2Ziji06IsIoct4tutVynVhLoVOTv301
cWIWUOmLutJBm8ta4bf86Yt19DwvhPhncIN+QE+nI/3D3PZUOoI2SN+jgt77++DO
5yhx6Fow6f+ZPJQmsKf9K/T3k40n/SG8W1oh8bdQWoyC19hee+jfSZXQfD7fPvH2
itjbK2CgwGX4OYdbDCCglbF1DF9/LQDO9+T5BZ88Q2J10LDQPSeoF72zo8pVT2Dd
q7uXXGD8vyk5iaqtCDJiOo/QcsXap9ehyBsVaPbQKaVHROlJ680AeQ8sQYgNWrxO
kQkCvv7qFO7PgTsYVM5EVRs98tgZUYj0mqkKOurEei6hVPPpQ85qAeujszb62UCX
PSKhIYMAnQRi9/niz+G/bvY3ixzaGFTEx7tgVk6vXUgfNAMxF2q3lZkBCSO1IVsq
pGxxNSMtqe0a7i++akhsDB9+1HZGt1n+SI+2QEHrY1NZ/upGCOkimR6sPVLN1S1r
AmJ9/dAHE3xvCyY2AGJLbqIhHhmGwkVmNQutLOuBXFlGs9Jr4i2lF8tNvzHdbL77
WjdAd5qRgNzAWcAmvMfXIRp8oBkTNVDNyAl8nvwciApuJ5Tu6EFT5GlyqXGEYGeI
7cp31m5yY0ovkLcmQR3tP9gKeoV35cUDZCKokVf3OafUcq7Ib6ttsr1M87aDjuLf
J1utwN/eUrtNH457vJiZhGDVloInHWAMbAlAC3u93AzSUs5bJvbc9nYpIIYhEfSv
HLPB4VSM/hRDuna8iPElFn/7+Wa8pw8g1ZJp1eDyQuetNhql5GQ9PMj/3smdwPOp
9qTRKfNccOi/Lmp+X6b15jox+QxZnzsw+QXBqB2FZGpxu7MDiuMIuvf13JClbXlq
X5t4Pmi31+kbsWZSpc81AC4dCrq5fprZ+TfiC9tG+r2iMvbQKAjHtFiKd5fKdOQM
DSTtrEb4TunryRB0/kVrmIdfg5azBepnkG19oYcsG25b7tvzpw2FnV3hOKloIjq5
ywjnLUweRmJ8vXDmTAxhcVATN+79y+XT2rTNBdPy9rpQgl1hCbo0LsP7mZNKM5/h
ENvBjHlBc31IR67rLruBa6Qrmf7G8LmSkEjYhuK0yNk9siwMefFkYz25FeEKv39X
DIgwQC3JoC3xM1/3eOMgMwlc/5gZtFKV2maIxtD7f3KbLDrP8HAV10xTZ678IgXR
AJYRCuwwdmuDUOeQqon7d3WDdl4FpwpX4/KMGLcGYrseaSserZ3XbHTmR+i9GGR4
6QTlVyuc9vsjf87lA5wWZA+xa59svf85oH6POyXDrIPu6vGv5VxHLa7USfn0AqAP
Svxhbz0BHn1kSWfN28ttN//4yV7ovv5we+2RWrvc16Ljuda2BIqKrCvvZdbOIBtP
FAsf8Jq3ioZewG+cL/QE5TkNAyO2dJPfHLQtQY5b5v+8pYMHwUnlJfIsI/Ybk3MG
8Lb0Ihx0e8p7cLuldHcr5c/+IDywukg2Zku39jaADoJ1QWngqz6mBYsI0F6LJbc5
+f4HLO83FOpyux1vXF6BCpc5JNaB1glRT4z+XmQsW+9YwD/iI6WjGA/hqU45L43v
F8IYiTIxVcxan+vOa97VWPPi0KUnh9sUBGKOZV/BgqDQzQBd1DEzy2z/7a5GCcoW
IwUkw9pN1KqWMdiq34UowPCANbntE7Vo0Qnv0WvOjXx716PcjDXvkBIzRJcDf974
C17iyymVE2K4aMCe7lH3Uu3UpOa2WXq2ptIn0XJhjmKU5tuMDTx3h6g32YAyyhVP
wH/XmqqfI6EaLGjF2Ma0yRhtI6oDJGhOJvfkTBwormXNRIo2Nme8njvr0RnXEoR5
7i2QzPNW1xA6KGHjcolkpd7W/cKvEH24gLarvt0RUup/6KcYo6bH+enbDicxIXZK
`protect END_PROTECTED
