`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eZEswf7uz/+HDs2YadZzRgCR8G50qEcKF43L8LhiRILyyV9PzjHG8mhaDx0+555H
ujvx1mrzlMeh68Q11pj1g3kg7dUPxMNcEsT6iwPjzEpRCNLhuDLO3AqfEoBXw6K0
LNwfK/AtA/zJhdIzDzckcfx+WtEAwgah/IVWZ8OgevC2uZ7YRQamLOd/9HIMGiTa
OT3a6Dx8TESL5FNJMT99CmGPAv0VjqSQWILSgTAmjsAribvg0YV+5XudGrltJ0ud
PP57wDQ0F5lLQCDgXUPpwwWDXN5x6WnsQpjBCvspcp0XJrt9qMbiIPB4Q+ej/fFu
cqb/SYn8dMQe8DfMQ9O45DR6fs1b7cm36rzHtnnm38JtQLeyhCsTSjsNV/p/odTK
YZbQyDhC8RNP7bL9HMKEa1dMFuYeuAXfiQ6yNeSB66hbt1BI/fProDDY2W8AeZJ0
1ds4LFYcFvt8h+RHYfyQ27qHIvsOTr/CubaY9gTBxe6k/IY0NtnGZRQRoC5o4bPG
QdIdGY4XS/dVV9o/jnsQcbKkqNYdPr1f7eGlkt+T6MMkf2gquEav2yEVUrE9C7np
oaIoskfTHNKxtHbKwa3YC4B38FGVQF3qOerelGAW0Plm81K7QFqP5jp2UJfQDqqJ
mpZ72K+R+34nP+aWPCAncNJoUpmmQ1GWp8KNlNYbMZlbJLvx+Yb3nPm2bk4HoZeu
vtDiBF4PEzUqh3QUl5cC+o27yeq1AM9H9iGDWxoeN/zcpc40j+XWYKMb8O3L9R/I
udb68bu8J/zHkfcKdcCxClQ66uxlnnIrwFhT48zLxgUXF+Eqk1YQmLrOU++Y2AE7
xzBMBajVoeojj9gJ7PeTmLgJbiBVEKrmAuGzxces8dqo9O1U3vcDDH6W3xYncs1f
q8FlQx2OmImKxY4kJ7fPkKb8IkZZAEGaMze6CD3oKLSv0wkkTAUK3MRNN4dwXHJU
882Rul0jfPr6j/9f4HEeyJQQIBPslsSSdt6k0PCgiXiLIzIPILaJE3bbYfTPCejk
v3rWw/bjBd7Hf8Rj76fElaCGyLl+BdMXPSZWmogJn5mPJ0jd1dIjSw8NY7Kj458f
qpQEKuWioai7fe7w1FnmysjhZi4WQCeH0ZgtOYG+RJoR/9K7mxM2xEToF4cjZFDI
5zn9LJHU2Vh/XlepZs9WZqUtpuW9A52s2JmrZGzxE+S5JRzpmQECby9H+roiGhzw
vMuAshdUsxMbSqROeqobHE534sUx1SrSOs/5Jr/e4u2U6fntPjgfov8QgBENIDD+
r5fJN53z/iUbJ/3XhdDX8coAhf3KxVDBUTP9kuhf4bzCTYG737cRnC+9FjQiWJAf
bNVj1tsxAebsyEM/xihp/ag5l1uoHCCYRRpX5oMRdd3/pWsqQ5LujwR7YDgAiRIz
kZmUBAUeLrpWXqQKvKkVnoGyNVVDh+oADd1vDQvbDtoxmPdiyTh6E03wKh6snbmz
kz9FwXaLts2aytgGHKP8Y/ytUhRF6NznD0oWTWJqMi89mzfe0xEAPuLW9iy/UbjE
k1W055qsAp9XrDn7pcwb7Pg59JKWR/2JRVTw8rv0bmtH0PwVTovvu4asSlCk+HhQ
oQQNLDK3Neqf0RlzjRFfBUoZPJfcSOfYJZhjRV4O4d3YSZKPRaJ7uaqEx7zfw/NQ
2wdQmwp+vatDh9AaAptRIDIl1p63Ynx0S4mgb9OksEQQZNZYOF2o4XYzVcrn8fE5
jKDSWsOYL+IBm+veyCGX1SQXFnIRpKaRfXB/O1VJLc2yVfuWTv2kPCwURNgQyT++
LM/C8dqi744qhG5QIgSRY3sVns9d0pfLyJ5GdxNyf46OGVvurJLfmtLT3Wagdq1H
s02chHfhQzxDi0pIZ9KZ9ieV3sy3bT9ulx6XZZyZQhL6EE/7TuHp0XCyKniE2LTG
/QHJDwao/7OVBE7UEZABsi1pqHG8TcLjS3Olu43av2AWbk2JyjZkVm8B9YE8pZo/
7g9LJWWPRo5x7Jo1swUYjcZJ/EOg8aWcFeYk1ZqMvXxWMSCPflVTkHKUQI7Nq479
9QFvTijuabhbbO2bMh5PuFOUtB4SKDmmyJb/VpzZcOrXVr6n34JIL+ZvXjmBM9Ql
pi76WxoNQw4yXKFxTyFDW895/H5f8JEKIP2h5HoxXjWIeM69f4ViNvqUIhGbaron
Ha0qXehr2TWtIbuahD7e9jxQAUmfieo2mi1lsqXbo6HuxJsOIBm1KnnAVz7lJdsW
lqhzZl0z0afFQ8xfTMQe7ht8MWMwn26pdLU8FJraBvo6cMnahYBEX3idzCNshCf0
rVtPWp5uUxY8o13hm5E4JZKhiZ+iDaYbU32AisL6il/0sUGYJCY3zDkiv+CdRonJ
gAgVEV1oytgbtU8b9+TxIzeEGHyO4Rft+yuc2oiJKBUGM8FKg8eMYFtzMUVwZVz7
1QyDh6A2fkfVSNFE/aUPNUJXigH47ZHE+GSxqk63MtLbex7pgPirI3bks1utGFH2
1OuZDGuqDyhbMI8IUpt60Hg0xBWfQhdxGrAX1+BqA/b4j5239R2638+pKPjw8R4c
pS0IZ0RcIAx8AdPJUU3cO01J04RpQFdFMQfUho07bsE+9yF9nOc5c2b19bJDAl5V
CFsIdmgHjNDLMuytZKCt9rMErMlEfKYIs+H6Q5cWf/JhLFJ2/lPk6zF79EbHnomk
Wkegt6zADh64Y9xZLVFQiOZHQ8eE5juHIzbYmjU9TE0u5Q2T7ztWUzCrtmoysQ8w
sOLFLhzzPl9ZDIDR3WEto9YAE/Y9EaJ31o4+Z5h6I5oz37kS1QAzkinrxJewQLJJ
NHKJEhxDos5Wfaw23qYcReJeuzhEsZBQysl3MKRX8McHQzdBAedCporPeNBraFlk
Dxqk6InAKJLfxGCiY0wyZ5f6knXhY96hhOD6QNN8LOXqMCS9EWrfgRTSkifOnHkc
kiq876Hhearo5wAgPu7ATVQXPGAss1LT4JhgPqbK+AL2kFQIilq8yTeK4/O9on8N
WgF5NIQ66p7puk4Jpu36Iqc4N1KE74cZjLcv316nftDf3jNAwfoNpYXcvXWi0Lf1
+tTIdEsq+bDG6xsbgfYp2xzC6McmaqzngfFVjnJNSLaraFDcPsMFq8YkOou/7Fix
wy4o4Wftz6SsuH53BH7Un9kIjUme9hsdjp4mxIP/r6vN4aDDw9puHdukO8K7OPDg
gCrb/ZHF6Uf9vRLTBL3KgBc0JHNkyvwGeUh/nC+xpZnAAfu0U69mQqiio8Po0yl6
H+RUSehQlZVMOfBIIdDcsP34DsL7BOtXrgugOh1JTSul2xg63SsmJbcEdsS7SuLh
07kFf5eIIfx+zmQoN+nTX2P+FShbxiCc8HEapvxk2ZRcldhdiqMsBUH/B5n7qR6f
PHOEgdTZndJyxKdaxYjNU4I3tmCGyoA2gYSLmUaeFzYeJogFr5yDCyBQtiAfm8uv
AgDBo29IoUKcmSjJuh4Tpxe+hyGDmdInePIdleZ4hbSS27XH7ybvC/jIhDqe5QOj
ydsa82Uh4BDtqYZ2/yrK34BQ/JrceMQ4n3LYWvwBloPa6nkm1ZrjyuB8GLPCvz8N
35EdpCmRDn7mQSA+tVQVeJROsBEPlrrNfra7DBrZtV7rDPHgBcU6kp9CPDZMFvvw
IENjCDEEGIv4xUo9rNqkdZ2hpr+iMnbotCVl1aBvWXfEDJ/8tqLqOPBEVa7Jea7Z
M+BtyxXh4kUFMG6hhd+WfnmplrF3Nh1JqmfIMTYaAWV2vscqtdxvvfBLj3Q0HOdq
SmbzkGisj+LMBD4MCBHc0376kGgP7F1WbUjYpPPkWZoiUXPBa51sZ5O0CTEvregY
v6aRngM8xUnv7k7YHyUjHpvQQLBmr/0gddivt44DuSG4952X0mLAxvT8BAagBihd
uWdT7OSTjQODIjj0+p3zPyeq64vBD1DkxdenZYYcqcRJd8GOxo6qwQgGRHe2osX3
qDBIwHWqjTGACW9isn57UHxS6s8SIph24BgQyfwCfoBf0/com9iK1yeXno4Oedom
9Co5QTvcjKVjWjsUipRatQYo2auD6gc8Ow07lv7LsIifx7TjSEVCdpxB1kzmeyNS
VHkKC40E3B0SaAca0YTK2DLtS/ksEUrzUgeiZR//BYJq0st204EVEiLYvhlzKSZu
8RDoyZqDD5Fa2SFgFjEDVgj2AGdjMo3E3ekuIjPzO25CRDnCbcLC+snkeANXhtTZ
BTL2vsHBLuaOLM8Ck+yBNmHgRa9CjxaKZts/11ox0oemVq24aicyVlwPHbFRivrg
1+sq7SkB8KIAI4pkxUOSll0OCvfwaIIS6a+nYKjy+WlP9Pk7q3AgtJMof1EEHoXc
EfUDyOLGuaiFIXk7FdqJVHd2IogiuPgLp8HKJW8EBGh+PTucr68Zom93/LfcYAhi
MP40/aimlKb3GvoGxK7YQ+0hysaRb3CI6KsUUBrkLywcNPWNqbLhHrSVn9WVpmS9
rwp+7hDY1tcxLwACwIbMCTMhRRiOOMaDL3x83A9a0+o8SbXR+BSm0hLXQ6u7OCAR
tz3skOyRGBQN6dl9NjorlqoFQxVXlS5kpOfaqmS6ky73aFT/WEnqCXSS/TFz7O/8
efc4NqrOO8LSZNpYi8gCP3qSVj7QH8hllKevm5bfUi9CbjpbgbP0v4PfG6VaQto6
gU1h/99wjiqOoiJfq4WGBiYk4r0a1IgAhiafILsvnTwFU3h6/9B396loVrGg1TRM
xs88twfgd8oEAbH5m9ZhTOEJRgzemX8/C2H0ZYePztUn3/njZn7UapQF1da0OW3E
GrwXin55dpOxdbO0+9hnxORRkdxp8ul4D712g0D2cKamaW2G8njduEUERpKJ+FlA
LNUU3hFu1Cz4aegv6fxndAQz8jSVGyx5bYJ1WPeEBS1wXlxqoXDCmRBQHFwut8vO
7NkmYMERl2DpXqJG7b8Nfm0UB60aBH458oNH4TJiE1AoMZ38S3jHyGmm0lWBIS6G
yAWM6rAZ3A5BgndqwLnE52TUfBKXuUN1V/ITCfDaTpS73tSt0ZU/6FCcMiCMzVpk
Bld5KezQYmsGYn8GlGU7aHAS/g4oglus8XDpmwxFuke4HTy9ZMHf3eofCjX+EnXT
i5l6ECaaSWtF0qvHSQ+y1YgVuowcWviwcZfoYy5PJ+nj60RWA/YhwNhZ9hXJJIP7
kDbsaYeBgDkcnd1DwumHoNAPzmz71W2uFW7LA13U5vKj3Ji4UBBCB65Xe6leHGPM
NdIBGRtwD2zP1E8flaIjF9US+v1b4EAsRm8hHikkV2o8HXBrFCdqxVCkYuXbhYn5
ht+2N2Wl9R4CJGmIhiiCQTqKLRVe7ifbu97+sBIFfYtgrqXwVkj4eER/jwsOi2LJ
UeE3qBju34TXsDM00i8XZWOGfAveblw64r1fJhR6mjgb81iRs55e95cHEjXAiMA9
9oBYG9fK3mZcFtDojy3q+mBAM6d5ljniPiW5pI7KQUvmi0T1qpTz227A4aaO007G
qIKK5r4lMmbOPuPse+eSNqTAzurXiO0QDMr00XM8tbQANhjDEbZmH+F+wvvU+9Ie
JMSsfCLtZqfEFx7dCG+HDNSEwYuOtgkTDXSpUgUX2xzg7L1zEj3UgN6NEbQgeocy
kBsJBS0Tgts1F1DOcIQ6pYmtiZbgD49afclvfLqyXfyHpN+mu68r5HhW/zCkuCmu
KDA5mjUtFMfSOAiQ73h1hpqSVC3Z42E44EPp45bLEu4KzdNbS31wsTF6vH3Y14Vv
6zysduU+j2C0PUNqPWjCkWunV8dU1Io7Gf8YiU+ka/MnREj4Kzah2SH928W/rCUi
SGCr1hvR5c1xWpzy2qzUPuijrUeL+Dfzf3Gy+7MB6vjkibJXYgR9A6KCa0h40/Tz
jaWF+l9MhVWQ96S02Fx45ZPwuWzM8zEmbE1h7Vz6mFLE7Y9MxgUpP4SW6BcVL/ZA
j1Ci3QNHpVX5QEfvdtFrUXkxSohUfUtu+5hsiw/3mUiUt+i/Q1pmrn2wJQwCKVbt
eB0liEUYgRpSriA97sGN5TU2QJCk60BXGuzdV7fDEG8=
`protect END_PROTECTED
