`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiD4uux5tlERO2eeGt0XxOY1+JAj6uYQ4wsO2i7yb4UNkinjYedUuWMmemsrYteC
pEi45KxOgVnYIQ39xK2WpfZEjcmazY/tuc0B3HRabWSOVsXaaqlbNEempARVLTb/
abnINgkA4QZWThYrIsCC3msLojCXj5OPEfJO9wzdqK3M4NwuJ3h2K8IhgqM9t90w
UIREHh1ORO4tDu0K56sEx9oCI4CrAc52uDXJnSzKtu9ELG8nCDJqWmuHAoX2WzF8
tTjHjUTsPBGlOGz67GOQRcaw1XttDrU2CxvgWX7Lll8GUCtbOohFoIe50HG3O+zE
v2c8qu+GTBIAirOelxa3dpI9P2FkTgIUVnuSH+p8bk6BpUB6xPgY6SH9tsCMzWXM
Ev9lieVn6xjCAPgC5AUl8j09QMo3+UMICrCGw4Iue2s/efQ5pwT+RwFFb8eiZrqj
XZAUHrNqGqSvU79ypd2zemwrC/rpYHt8DYCZaNLvJFvov7VLKeW+dtAEZ0zObhQg
dAknM7rRe1ORgx/AfuQknEYyt/jAxnTz5PNJy3KD9j9TaObT12BGhltMbsVF++cM
xCFU1VH6h++F3ANojVxIKuYGlYkvtCgdPBEJ7sjV9GW54BlgmVPTgLLUBPHawVqI
+M5NC6a/AFdjbCcJKv405Ti14wssWKzKL1/BTV8Y3ZyWngDKb5naVFmm2pA6oIQt
VYTX0Sf335PYvcMRMBeiyEpTTrJoLSvUGrz7GjW8D0/YwsuNDRWz3PxwZe6E8PC5
ysuMaVwJ5M7enUVjQ53SixnVtM6/AYMzMJbgV0uIS1DylSyYcvHZvnV3gMIwev49
tai7JgO0kdrc2Z0adgdetJW8m3XHyhUzorTh7RIZBwaLWuaxwwtN2bK7ci8cMCwY
qT/1QoJnmIa7avGqqb17oxqO2FJgnpRw4bDFH9hNPUcuQPEwR9PQeroZ0OqL3HGc
lJhSGYTI6VqH4rsmb+qSbl2ytVWzr7n7R6ClCdZZRYlOWsReE0FNqn5pE0rNei0n
wsTazZFUhlCB1L93M26W8FnDScadE077Uos4rg5sKDrip935lDJIYj3xGibWkQEL
fVscT88OwndGfZV0VC+FlGiv9x58H/EcX7A+feZfA6ik6sUJC1HoY3GpgkcgyHC8
QqUcfpeAoEJ4ijjeRli/ygqwESrKjzk3M3gBIjLZ9qD8NSLaQIUEfyXfirnGIc4x
JXfAQYz4UdmTK7QN24FWrgvl3G/ZoLa/LrqtLl2wUyRwj4++CMSmH1k3cSYJsvRT
xl0GkzF1OKFVK0g0ZwEK11CPc59CGr/+DkpIUTRL8KBtxLw4YKbFZwrhhgCejz3l
lqe9TOCgKBoWjcgpy8Cay0sCH3PZWReMi2EdY9X3KTdQabcTb/9zaoFe23XL5kIH
RM2ZlJKH22XbrXuT3bpLlPJy/jo/cbhPXItDd8Aea6lucf792yyvJ5Nh4kKbCPiY
89utS9kHcktRv+xtdwe1dqzX2rwTSLYcWzydEr90X+P4X8/r2NtyIamKFHY7pHA9
uhVnFS+Myi1fYikcdsBhOQw8sFps5yOMNnACg2IHRxhRanhlLgZ10CIV9+cvhLer
HKEWehFWkYFC2sfec8NQWoeKW5/klLkBGf2G6fVjxW4cIHYeguiygL8kFUunh7Vg
rOJlP7p8XNWawYzP6XTplbcfcLYX328bRIfF67wQcaNkraI7odPP0BGQZBkQNZ/W
+OQ1AdL/gLKhIIxkiOhvdbwaTnHTD3fQFdGrgHelzh1wHlEofT6w+lGtGrpMhcCT
QBtejEylFMXUMAZ/S+NGZFIfLgQHqE85DBeKbwETV8QQmAXyPY+buWw8osaQkFuS
7lM+uTul/8cI0zySbP/Ykqda9GpyU7Fw6DFSPUskGPANtPZsNZ87P+KPp4NHa3QZ
s4HsXvaesahkqoijI+roFV1j2K2gcSmqAUIbgQ1h1JU5iA/s3McABZxVkEKxo50X
b7YR4vUM48+rB3bPFyz0ah6k0I9NQHlbrj7PjjTqW+oyukCGGoyOuTFqkfvuoM+2
wUZj4fHgsphuaBD0dIsCJAN8lwXwj0M5DCccJYhT1Yu5uTAVLGfpRT1wuNF9uCjG
sHsqN4Z5zwJ4Tnnmz3jUfahOTeAuOT8CY7VE01zsWIn0GYBGZzuxMqNuPZfn4G03
XjHSH8i36TAhg05w9yTPW/6VdqWKUmKcZV5AYybBziBjDtzvP3yPfdCxNnjEZwfb
Aa3h7NOS5J2xIrLe1rFAqPrFgWuFqwyvE3ndyg/1R89chnqMriDOi9+1AOkeBCk4
2l0tEUjtqqkx+sq426h0+inagF3c2Tk6V/oCUO0w6pF7udL6MTi3O2PeqVP0w5H0
WLNm4hu70T+Ma9w0IyRaLLdQk00XUvDXA6quLK9Ma8vICbv7RiMkmWzu0LkT7F6b
1DWoaqYrzjGjf1qw39s8Om5Ynzi0QNcl5MvWXLl0L44+jPLrx50ZfvURd2yYTblq
47Ljf5X1FYYAi9YY88HHkbYgYDTvWgKLZF3Rl3H1L8oV9iSkPN8iVxHxgEPJa8bc
VAYX02+x7l+u3lox3y9NB54oY618jgPfXiW0flCZGQhaHVSR/lk1zDwdYMA5LK8R
/DhqSe22IsyRK1qnIDHwauhFjp5Fdvn07XKmzBX7IWjVaF0l1HfDHX2G20N1uiuK
7VRtvHB7NT0Rj8/j/fL/Epz82fW47+rVtVVoKrcFE+p1T0SkD6tPiW4Yg8r2euEw
vS57H3ezT7hKMyei45KaXv6gBRrn/hHvt2H3U4Dfp7VuMi00Bp+Lx2RYQGtNVslV
fsXtDuLLYizk5kgPiNdFVeIcsM+6eIi/nqWbLqIwxXuZZ+o8YGivto3G6115+EdR
FK5yt5JhuHqRGIlICUHU81M8fywvkIYBvxXDtKOPuQ7zMH/KCnkGN25891Yr8IsK
L2H/Yoh42xVjQLeuoBUQ6NO3BYtvTmodQ2+/6thQXoccLK6gnqSvkQUg4eMI6MN2
mkaSxASy2ugzsoy1Iv8isn9/V58Go6Pj2bumZBdfKtcWlCr9kHwnGIildr4bKlUG
abGkcUOAY6fITrg6zj+BQAz2gu8szP40s4zPYZmg4h3+KPTsnDZwDAzG489OsIya
/pyVEU8yDBrDbMxSpr+IP8PwEWPObDz0R8+5KNHsKBvG6RG4PcM5uI4SO4vGZGaL
affrrc8VO2hVWH6G8biidl2UiqQVcLbqcNCrq+9edPLOO6oJQTm+nlc65uo/moC9
TJzx5GIye1UQJnwSz8Ewe8mQFQSjFvDHmbXFDi469ekaVmyoRaCtQKQfC7Dcx95V
F9ronGOzi3/DmFX5PJpJ+2KIkmyUiv796JunlTOm5Eir+OzRfNN3PR1Awif81YJq
Z2+gP2kr4f4Ruow/8uydGeipZa+9wYR6gqiqBAIYpRzX6RxTJsPxoB6U4yhjbvDg
H8FJhDdd+cRUp1Md5IXqb6lZwK0Axl+WwY0yGfNDAV4vwOeHX6ATF3TJMLzfikfx
LGlipzHg5QJqqw/ggDQLDA8qFUcJDKVjdwJ/5gtacSbEe0Bc2PA0jGjFxCWuEe1V
n759bAJhg8n/amLupHYGsZpMojl5saNPAnEd0WRyLvNvTg2pkyCnmXvdh75KJUsa
gnanQN+Y7XLT/Tz902vzQWueBENxVxfOcaKD0Qdz0xB5DuU82MBFmQOyv+X5tz+I
7EdikRCjzqmDKurHxcgrM7+ksHikOfc1VZqtLfxIT+zI5CqxIbiitjFiG6L4A3L+
Sbs0TwvsQjxoINTwXlD6uyXvXAFZa4enJPKqN/cbMyWAK62DsE43fy3w02kRLTrY
tz+uyZtdw6M8cSUJmH0Tn/KWxXLJBu17Ng1yqxujfWt6tFxHxlW0paDxIXFFOPfN
3i5m+Oj71SJiPhpXkoTuxrGR2pKIeimkZPNVCJqGmsUNxjUyInSlMq58d2UP4oi9
S3/2+WEARhgShli7qJHVQAR+C2rPGqKPOAiLO+qHvLK5nkS+RaYY1mfgRb/r8zdQ
vQfbfhWINrV0Y4kXBD5imapqV+6vNOw20g9f5AJFKYGGhcC5ILgWaUx1p/2g68Ed
zCGfAEYa0kYBCH3XJlJh5WhJYFMlayGIPB1+W4HsSGXmLuzMUqBWp009ElNVRImE
8uBs0CBSVAq0Lhikh82cBnzH3mWjnMLCwNPE95PdM9wBz8kcYsn53R+GaYq82rT7
pdVCcgB/1pfkDCegO4MreLJFljcOhST2MB0isx/s9TY9Y1fjHGyesrNqCS5mLRog
EI8i666oSz3uwgdpapVCO5jM+ge3hqT4r3w7MYreKLoztwn7NC7L0CH1gwAvAvaj
FeigMjeiMoPamDb0yoS9aYfTE1o3AHPr6Iu9Y4ISCwFJwDo4sUyTVe6TstKwOlw7
jLPMhj74LL6niDHuCFAQ3PJevY1MFcXto7pesiLWztPCRe+LDaI0h/qCqY7WdBh7
oyid/xl+fxs0hYeXznbSutqM3GWQ3VmI4CRzyZO5mD1DJ4xWLvTKKz++wutIOV2W
JHoYe/1+Alb+tsY9YCf1NxfIqB7HzUUOQSSg9jKtcsC10o94hYCHsHwlPfgrv2mW
hnvffgkF3FmW309xq/JAFzAK5QC0DaIPoiwsuPblEdkk3nnlYkYp2WJBYva0BoVN
VzYdRztfUnx8H+bVsVmdMbLyCgJcRPjB9otNnGS+LuhbSsSOtgFJ6PhMlr6wDjdC
+48yTeaPBiib+LAd1QlQRxQ58N4vEoNQZZiJRKj39c55T4/UQ+gYEpvz9erbgpdd
JWUMs7w8EA6/aSPMbuteYgguL2Rw0mtjT8rHp3/s6O4D6inxyMoneidCplvkzK63
n1lRE/TGJ7LwRzz8kdH3fvmeHWtoHnBb4Lp1ZkXb77qyHf9N1ptV8kQaZT+QNymk
SQMbaT6nO49kvPxLVC8fkE+MuwfwCX+v0p4mST8mXrj6Uuzwa+vZQEnsI1Lna6ES
n1gCLL3Fq27CyCz758ZHmqx5GVapEvilaZ/xklIlChvkx0PLHXnko83aVmfiz5lv
OQmDIAGCEUu5WsTTzXCWX8oynlfrZC0bUBk7X30RLIoFi96rwiVNqrAWW+7R598x
ed1PYJYAfFXWip7Kt2MGEzyglmAukG+0otL224W05WT/ROBToXsqD4A6Eyl7I4aA
xYAeRxaOGGIQwvDj40E9sDaIujfGjauzGZrPTLM92mjKF/Z05zestJi+Jk+i7UG1
hXzBoUpmFg/1YLJHWxTEtzuHQRQnG3jTYm6r5W+8hupUHRgpAg7l86nGGeJTZ7AH
4kvh6uxdmBPohxO+HVEKPpVO8Bum2ddOxmnpIW7nsoq1DVGGTA3CRsciFy3rxYzk
rqxhLR+hud3Yn3VscRFDxIF4KONMBhQu6PPbzQ63iT2oOGqAJQdz84N34HiGjHI/
KkzGL68Zu6bYI93u/uo2rNhuFpiVkEnM9qzF8JiUDdq6lfEjBojMTUuV3Rd/6mNE
/8l09unMlqloTFh1TXrdaxtM6YWgJBWpH8npUX/tVkziID22BbBGBof/Zv3Q/WFf
B9+SIu5/qy1z57eVSmV7Ka8DeDIxuKdIjETz0FvQHWATxZynNwSBchKkKHQ57hA+
kR71xQcZ+Tn2/yfUMFmf9/DVP7jZxweb2yibp9f9JDt5ZcUt1lKvYeH1UX9g48km
T3VUAvNoPHaLghUzZ6QtOLL/JkPx+e54TA7edmKoBvZ4WjVPxC/urgFdgkBDIPz9
OGJeVzcrM45sHXMIp3YM+61SXJtzhWY/yU4396YRoi5BXXydf/hoE6S59PZn+NJn
upjHo0tsrIVIaBGsWl0zcyEDMGga+kdEzgskB9pppM/VsEAuHMTd/AigvE/Gxob7
uwZmpgjVs06IqsE8WO+SVeJYkWUkLrz1Go2b+RM1o8iwmTEs229uvGc4qbdGfX0H
cgpADdM2NMO6eMGbrft68mIt74/iaAfX2yXNxLP8/3qboNJytWPQOPkuzgPX5lck
5eJAquS6E8UcEfoyewzKb6v/X3P/9sW9MDuCyCc1pChqJirEMEBVveTuSI3IIdfK
jP960POFL3NnUy0sIFsbJMn/ZZhZPJY7bXrMwI/YXM47hWm5nTf8HZ5WXBRJ0YdT
voaCwC+YvZyhNqgmmKjPULYw5JCnDfw9EiRxpMZNr8CeQbJK8ZKcUcjHCcVmwv18
XpyP2M8kpShQKSx1gOAZQakZAbOMUGVIdOF/RYYg1upEJRJ6rrgOkHUsBsKD6tGU
tLDnUg/m3byE90fn0YS8Cb/QlyAWM930GE5xH+n6GveRsrCmmRoze6onx2TttwY7
2nnb0PshOlEXS9n2+SWSs3KT0fasbNo6CN5TGIu8T00h45MgUPYQiEmQiLw0WBlW
xhh3vRnA5BkkN1p7h1fzIkeNv7z51F7kEnbz5LLDI2kcg4gIXt4QkRwRWSp+glkC
K77vshzSm1kUiSYaTE/iq3UtTFD6cZ3CaKY5hyqImLi3erXMMy3VEGRgNGkgxcEv
0in1lofN8Ytty9ynk4cU77j/yyfKfBgYRBwh5ntIA9ZneDVtpxuwF6gG/F/m+dD9
U2uu6M793ijDtdKiifdLg86PWMlApDbda0yyfsyLtJ+9Znh2xoDskaiSrhwW9EJg
nxClsnsvOCYTHBvibjkZa2rG22F/O89GYDaowbnicfbuwu4zAE7O79XxJosFr/Qr
lpiC+qWWiBNtdCmLAp4WDg8fQ9/ndYYaVnUNdkfkeINfQIi6zF9qQU2OkadN9ubN
dL2Ps+vqiOeBvJvBpPimXNclxyCNiVjKv1m+rR2GeQIHsuJUCHEuKjH0pDJt0jhp
F6EQJKZxtKuKQEZlGb1kXrSjuoMUCuc2s+QNAnkhAb2odc+RC5ALfATnX0dSKJyw
iYLgB4vaZQFnRy8NT7Pbdo+jM8Ggc/IjUmh8B4YededlmKFts4Liq/K0DkBn/v6j
nUhkNR9UaufHOnUIX1INr77dq4YLH3m4u9zM9TyuJRc7WdrdLtOifTKfcmHFzkJT
oc/CSuHMjLd5e1EiHDt/H2wdcPvDfqe2WLkDM9GDrg3vjOBHCGQBTjmef5aw1Cmn
1bSzRmzdMn+5sjoAekACMpnYypnZb54dk2JIlFqRl+LivFXIewM37he5meAjKvao
bTATP2ffUJ/F2t5yV4kowFXuSyHT7rq9KC7Jl1zqFyYVX+IIf3+RcXfT8i/QNLvi
SqdcUtQh+/XQVQYYLkhB53T5IxlqDWPFyeYpYTdQfxnRcYDzSfWDFkEoLMUGiLyr
7xzKVLYPNbA0YCjGVq4M4MCnnE5xnfvoJ0BVYmsaCE5+OaUzm7bJaJYYnnfpy46G
VtsJz2X/wrp9HBp1Seawc5349+7zNGrzKRCPD6dEOSyRCJjXT3dd/MDU9WWHBPh4
h192Po3ku9D8mqUioMymLkxctQXxixXs5VgaUYEbZfZiTlswCtNFTTgPFcyqqjOG
lWCykOTvW5/MD8xHW3YGERPs9W/N43zKTf3LvJNKpBtAxn1vfgneUs/RvZ2lXdXL
L+dvKxu4NVEmEQvODWOvSvgD3//iGD6TLgDyrLSwZcyiPrZcjSLgWidRyWDxNVXS
QbXmRklgX5w/OnQrB/+MZhAO1FW1CuKazS9ehWcF4SjSk8UEDnkMR6KsiBxsKrdj
`protect END_PROTECTED
