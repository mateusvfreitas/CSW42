`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v4WtTqgGryqq1mtrGGbM+2m8rr+28vWOx9PT2FyELwlPx6J79W6Rx1iVwx1F83Pu
vchB/5rsi3GIelAfl/eB1S5wysDhh8cngcPrDLJNIMcRiso0Mx+QbDUmjY4tvI1L
ZVDdDz0qqj/shVwpJ0E0sTqXX5GSmRPsxM99LhIan5CrbpeST4VLj4Ayxa4v/58q
xQJXM+sGv34bx8j/BA/POQGrWG0Hwbxum03UBxDtuf/3FXPoMSn/YS+E5bV0smEt
UYREXrR0PBzCJoYL1E6ZBkEJajqg8YqRbGiMZ9c4ceWytXCjeHtLRON6gy6B0A8k
peEcFpI12wWqPvNpcJAQdpMhRi85jGs1mHaxVhZpVkTSK0Un1lHafKrDQFC41+jX
Gru4OGDo93iC0GqeYgCGmFJAW/3mecCOaacvW6Tid8XCV48VoJ7RQcKNlHCvFWbd
T2T3WuQ/0lxRV9h1lnIE0gRH2nE8oDsdbY03lUvsL1jYQL28yNXzvi9/A2xVL32L
wwNmDGAPpGrGYofgmPoNzxgs+lEOaY3DHhirEtpqeVcnVxwuneenJls7j86WKQLC
NJyMzZcZEbcTkkgG7Vf2E+UTjhRdiO4VZ3/BYue2g+WgTrk8YJKoV9BSBWVPD4wA
/pNmCL05me2J+UhvjOLzCX2dWtuR1sY+Uz8GxhpzbiDSnpLbJ0f+6/okt1MydjQU
ot0ZW2mJq5mrn53B6PmB/ZIxywdk+U/bzDRGwjAVysY=
`protect END_PROTECTED
