`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G93Xk1vsYQfHxN7TPPzYz8DjOCBnxiHMpU5mTmlDtZuBJTf+wRBdb6XKvPzb//zZ
2xU/wzfgtIDW/UVuaLi0ulAkZKMLH3e9mY9zlOqK4qgBnS71jZHqQsh3Wo5lOLMX
YiYZSTLhQqnGtPZSWyC4pJI9uyVS4cEa+zfTHSulIgWk62ZDnhMDcBmFOwhcfHHu
elGnKSBJjg6Q8nAIEqG31U5omO46CAZfIGCLkyY8rpnVCWZeQtEuRYomT8IGSTPs
CPJHUxjhVeK12CqoVBBdgSeDsW+Y3GunB0hD7RYy5Mo6cUwRocXWcka9TMO3uM2f
ntD2EujISOhlXNJAhG6xX6NsjRGBNdbpTsPrmLmtmrKztTu6LXfueC6LvmexEyg0
Gl+/CFo6iz/iEFq0N9wUlpHsbYYEY+P4g7EMV+RUffPajlDqrDr6k3uhr3BTre0E
GNkORe3wOPT8SUCO2cex0UMWDPiCWMqJ8imdgGxnn524FN4XHHcP4zjLdkyjUVve
Qot8XL/Lxe/wgrfmJ1Z0mhZ4EuDHfqJSWLDfpQ3jYVo3s0OMOgwE4lmvArblBD9V
rJAU/36vgpsCkvkkLueu7dl09/7Q6kTpXXmfzCnvuxh4kD+dSUWRp3U7Ji80OYs1
RSoyMvP+RqOqVnmZd2CAUu8xRgTtq8DZphkzSsrGZZjuxcMTcKEBngyelYyUWnqA
H+ih5OnY8paV+24Ehcv2uh3yzWkUBB0xgn2q52NZZV3SWEsBGJh3XNISZJEcEsO3
93uwVTJ44tRTxRunOEZjWONYXbdB1eXp+iCRZFO9SNA33WfzWp1na3Ic24pJX9Pr
iRu+vh04lF6B8efVXtIJG2bGplBqa3v3FAgX5kEErrFd5aII1RgFbNZ9QqUKi3qS
HiTOkL6NBUQrywwxyX1r7Yu/sY600G96ctMy+mLA+x7LfDfxXDjx2/3K1InnXgA+
e974hCWUjWvCflzgLK8J68Rbgj3Obgs0JK7u93BPQwTb7G1N0v9TEpWVtWVmbB+v
oL3b2h9c0C8H3k9+h5oj1Rzi0Eo5Hwqvlxuz5+3JMXFgD6p/gulNlJBsAfQL3YOV
GP5J1DXe8M+9/GEQpn3GfU284I4xRL6tigIMZ6HNKAKFn/tKOjiZKBGRmoCDpQXz
M3zFYWuJS7J63Xl4PAFeaJY9Gew3AlYDEG4xY08lRjxpIyPRxaBXeGF3vC+BGWwB
sNshRJNacY3i4q3P+muIjHuSOrHESQpY2HmdFX2n3TPJcfIpabsV5wX77TCTNCGb
QAPBciQZxKQyz5sab5n2gXz86xDrYeAp2nWQCCJSuygtW5vRJWhHLF3CpF+WcEuo
/O4aH/1mXyyvufcwHVh2ExGJT6krBqztZa4j+KOu6v48MB3/82jJrgKQUmVfeDuR
SaU5CE31TeCxBjYzdd1WnM8UpaCuFJIaQ+CbZ5Xf2Q8Q/MGmv2SZeQSL0VGjP+vP
DBJsh1zDK96mye8L44joVPfUpkVeONPCL30diZdHVbytRqGCpOqZYMZdO1G4kCk9
jr0ageR2q6hV0aL/IHlP2tk015cUGu9Nk+s1Oadj813zrX6W5BLD2pDKKvnGptgq
Cv6vHNmOQ/C1zebVU93Tf3RxZTnBkH8uGnb7TKVPXuCzRu9fK9UuHUbuLGAQ7cIp
aiBCnL7WX694TJ5MseArfgujrXxmWw+blFGRwmS3rAsclqO3tGBt85r1pzqbMeJx
blsFcjf1iSOmMNPRiBb8vhmITIGGpfUNaX5PDDXFmbiRMIpyCxBnN/hm495kfmbI
HKrZjga6hsavj3Qp+B4ChfryZFELM2Z4ZFkwxTwbb6eNYi029Sqlz+l6MrNET1EP
7MzOOgL/IFqwP2AX5txWNlUrsKpbyDSWu7Gj9gHWHtOsW2yCk5anKpa3h10rG4Dl
+1tRGi+uP9y4btGZKCA9NPRG/EtQ/6JYtakVTbI4vheHh2tJ3oIGdku980cFDhCg
SVe6M7X3UShjJT1kgi196JKBcV1Kg8yypTKRCdxiBOF1p446am53QMQwZQO3QNtZ
mW6OkQXEAw8A2N8GPkaXog0I4IBmLpWj002mcPWcRdk8psx4mW/C7xYaH0Rg15rk
ekbaPv9/iTzc1mxaZG5fLJObyVWLONfiRiAB7sm93p7i4+irrfQdPacaiMs2tn1n
EyBEUe+nZgQYA2nYc2GzeAU9yjNIwnbyg62aI79kLK64rZmLVb9Ypdh8PDg1iqus
7Fl3PT1mIJRe6zYE/se3JQ==
`protect END_PROTECTED
