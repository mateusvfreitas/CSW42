`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DnvB9cVjSCfZcGOqdRCMEe5xjl2hBf583YVQEJFrcnUOwI43wOy5KeaVVUGpfi3B
AdXqnR1y7PpZZOBSLVRFhfQoqLWROIYIeaPD/dQOsQJ/wq9xeXzR/jmHPSBaLhhz
nxP914WkOz/+UZnoxa0Q561RvJF520yUIXyPMBO1Rj73Oa+czsEazlBNQQViT+Mr
Ds7sRP6mNBlpw6WlggSClSDbjylrkmbtxoI3aeL2vdo3JUTsY2dvDe9ioJ6CMeh0
dGHc4KsST8dcupQKRG3gU8gp4MlGomaT46HHgb7V/PQdfbpOQOdA1c5VqL08q59r
ENRDuCoLD5wF2mTNql2OE8+cpy8cDdCGy4Qf+pOPWXyp3dBoLsIozDz3DVK9g6YC
5i2epW0Aj0cWwnAT/k35GCGRqDd6tZiQGI30le+Mvv87Y/PKy9p5q6X+wK68DNwc
0voPdwi+dVmO3vH4keJ50h2Lcn6VfxOA4HM3kgHVl/OXJ8RuW+vnn/Qbn4P7mINj
klm/ouBpa6urYRfDR2tpI0ySSPs0c4YeDMAsdvZph9CMyLCPvwZgFUav6533uLvZ
TncNHbDSPHhytfusGF1nPYqxWNk4TSTBPH8Sn3sSeBmqogmqGrzGJ6uugWSFpw3j
bkL3JhaL2SIXBGv9jF+amGGRoYPVbzOXAamBMgr54a3gzBGhDn/V2VTAlciViADV
YVUalRwxRwjK+xoJKY3Bxc6akq9sBKHy+l0SuTZtnI+1ritI3Z2ibOzm6L6k0lZP
MZTALQA5VofBxkcr9OHi083IgtSOFbvqJ+5e5oufEcsSP6HI7NvjjBGZ3Ur3O576
PzqjDQcCtRuKDoisy4vGambZy19HlgF3a1OZCpHkHJnRIxfy8RHOswMaLoEsBOws
1J7DkPzf9a2WJlABguJK98p1s2kZO0AdOY2NiGeu9l3GbOCjGoRVnTFgF5SQHE0M
6CfKhtM5F8yrDUD30arOSjYvNlhjNnJNPpcJe2GAdi6HhgYtVF4CBNuZX8N7w1Mo
+5M7fhNrnLPxdJQRcpm5ZaTsHaDreAhBOYrOkFtjelo3oDu05pCcvuZS2bs/sz8h
uyff8ABs2Gl6gNa6ymJvftaN7+r0z1Wbtlkq4/eSg6h1ib0eM2SjyM94pPVPQQhX
eQ032rG6lOE5fnqBYcBQjoixzKblwqJ0s9dHki/NO12lAYGPzlZVWSX4qONJZ47N
KzppiWxSQ6rHdipeszluCDcdxeD0T/ZXVGYbCatCnrzXwOuWWf+IN/immywlimhm
SDT+5gGfUae4vRiXNx81a4VLhuUN/xkt70y8EffgjD1nW4z3U8XemjSKIHeu48NC
Fek6Ofhm8gWFhDeVnhn9OUZmOGCyR1hljS268fThnbdxahONPpOzHQjyDpeGf/AE
J5TqE02B+7GhWlUFDyyLykp+IgtGWG/MRkXerHfcLv99mvP34QrbTal5Kw7s6EWI
51i9Auh9gKghqNo/8i4vGPr8Z1i7B6yWWgZf0FYcDVwUxhTUD1pnep12kJDSyiOS
TAlw2VLlgcVc+sUjohdQyzg5WJ3v+PB5g6dARQ/PxFohdNSbieI76xu8zeC4kFmS
ym2YNK+O5TaKtmfd2AOa7FjxdfoEyuWhLDN8W8LHfYK0k6POyXp/cTm7YnOaBsvJ
8Wzr9GN8U7+Mji5325suT+65JxF8eW1u9WkDs3VSbnHIBpU/Fv0jVYUEqzLmQnp3
phs8RYqVXCY1p/0HHRRfx+4P5c737JTOp4dFTBaVGvwfgN0KFOS2iH0SZ2esK+8m
hfHY0j2/yMRkypNw30096CiOrXXEUIGiRqKLeNlo5EajlTy72bqC5PxaJZyC2SYn
9vnBwRYtLK2pZI1wjhI7YTNBavF2xhd7NkMO50+16YNDVqGZfjWOlWPk+wfbKufo
rQOEw4kSIv3KkIWGaMkOMqKChRhVTiCcLnZeOOFbonvTbkRM8G0EhDEdxdCXLJ/5
n9Yee5snXBW6cW1tqToKxEyi75ZE4RWW6c69LsDhHlzYm8bV0130r2EDjJTqFYWu
Q/Za5pDgeCzh5A/rFco0W7B96ywgHzsi5RWeNhNfTuObIvQvFXGCvohTeK32uWR9
pOjiyOamKBjvmiUfubHN3YVseaarzON0DQal7eE3vRuOoCh3QY/5uNUkM02EYMKc
mjvNaSefyrsB0gNgLRGxI8MKT58gUICyNtGhphPi6bf9XcL6BOUukzpt9YA2ZOf8
nHdYGU65pgFT5C1wqUWh3mxFZGfM9jlt2aP9y99ilVzJe1MNQmn/qqwOtC0cTu+Q
eQGwE/ow0LLcpkGCXRJtHqPHyLyW6ylENBoEoIzyOvT1g/Qp9PKD2CFGSI5Alhr7
C5h7Hh46V4g1E+fNwwYFf0sbg0kRkVxbYWngBR4sIEupetMRR1XSGB7pwxyaa7VB
ZFyy9RviXFxOqF/9u66hgpQ1fEhM43tEXkfsOBw6wTGrEGAb6s+kRJj20iCJEOSk
J+JiWqFWG4viHTdUkKGQd2oZc0jAqU3GW7Q22fnd/uSTD7vEpBPZrT1O7a26nLMf
JLEWkd0GKh1cZ+Dg0EcPHfvDAv1B0FjaebmMGQ1hCkRFvhaHOiZDvq8Pwh9iv4lO
IKWC+yrMqV6eN2PiiGay5SSK3lL2iwLZ0tjWaUCzM9/pcyXiBDLHXoyl/lo5Lj8n
tWm74Wk2Z2UMAoPNXV/g0rZtuJJYa3B5ucQ8HKYfQUyjUapVktTjr2UabYKK3Zhe
LeiRFq8Kd+ynQbA2LWk4qdWngk+q2aAKQSOkx/Xrj1X28W6MvwFWpF79dZONr1tc
XZbzNPp1f7aSeyhTbGJNVueMoTW6VS2GqmtFUlm9XVbbHxaD6qekqshLUBX1nlXq
HGHGPKLT8oL68ZX7+moU1MKiuOwW2xaDjzM1Blck+Vn39quwHezSXouirfp44eCX
+Mkp9Q3Akqgw0J1Z3ROSOrhfI5nXk6FBnddPIvb9hVrQMRyFfp7C+vO2luuRNzdv
RvDjE7dXkWOjbJXWqZjPPJpPEQnaj25AE5nigwGxLPEX8cvgowm+HhRE6ehk6ufq
5FotGVT4IVp7jXXH523tJJyf5wsLxLIdgYyu5XtmvQFTFxM6WQQE/y6FgCO8yAgV
kx0UUMr2UWb1L/akWzoDhRvdqsFE9eBTrRUo3uBe25Tgytmw8ZfbW6NzirVbaS5N
OSj62r3AdrMllJeT9rXmOhwRhQSWWqpWZcIZWjTl21KahaXIOhtsPjUvqACWrR8b
ABPb/Tp7IJDI7X+q+d5ABXyFm8/z8ZmR9RBg5Yb1TQIThLwjKOPfIW2bNyg/q0fn
6fuNYFI7OuPKjY9DPYZyn8Xb5zfv3Q6PvtkNsEn1PeQywfd2zs2wGh0a6ZkVN3Or
S5s0hRlNFMoycRk0wcpLSE4VIGslgpjcr22zxT4wVq0OkrcV2ZloYAzEjRDaCdwl
PocLApwE69BcNWn1oILtsrqSw1+NlcUgwU5poIlVDN9N43t0n9nIuykhlFIDLFk0
iBjGBjlK3Dy+S8/RTntVE8rXRsU8m1iDyiwbkS7WJm7/9TWNhpdxz19BjCJnoA9o
mr4aE3dA9Rx1dORnxBfe6zIYmaoqxU6OJ2+5Ol5UMTWS+HJbnL5/jhK/sJJVBlbu
17N2/hWynEkTkpHITt7hRMIne33822vOtqiLRvopRQDJoMb465hoVN6b4wp1WKB4
gVOku/NawMdctJp27za3s4+kSmuhJpTVJ+4wmVjBZlC/5vSO2sA5IxOYr5DzjKqB
g/eJGn9mzpqG9QI8fW5LqfYavt0ypIYJwog7PrZ90H4XD8VLnnA6tsKAxOojXRWQ
ShffQlWK2gfwNp4lSLWAsIp54a5e+98Qi4aNV4l/DAG0Posqok64eFnaK2qG8hyf
M+2ID4OBjC3NaqZPSgA30X4WmCQOYqs4LUSLUjC+naXUh2Q1tguy4ojePVdgOOKj
S0wGaHXM18Ty9v7KTPlUz/0wMvrmmvEGifBM01GYNGydgaI02XN6G555n2oRLKIh
bONdpqe5SsH+HKmzs3vmJ0zUX7Gg/CSmtCp5kzn9tD21ROLy3iElcfWQArlPAyvy
vVnjO/TV92kpzjblLu/UC453DtaylPad3ARSb8sazGIq85Dr6VQk4jxKkHkV+oOr
FebidhdKQBkN2zObcG+AG6xqqkEFYRqqHc0hUNAwC/5cOgxDFBiF8S7LD2Cg7zjg
dheP5UWEPlOyeQIy+PfD8hsIqs9rFaT1U3RJMFicCFIjIuVgDO7uGwh2TEXZMhm0
V713bvyxDIp7jTWDMtz3HParxg3B98wqZlJRIwz/fSequXo1EiRAHSAY9G++8LWo
4ckgJPhNI0PvU3i4Gd1ixLAXt0oiAfoLo4qlARdFfCRkGawc85SupVBSJkwmCGga
vvF9iipQq9ijpGJ8de9yuD+gV3B1NvcXtcpDOo1gvOUahJBvnHRJvKROdO6Lrk0n
8ZLr84iz6XgMcgwh9cUdakHNRVtuqzMuFZI4Q9vH/p/W3KkkT81wm3Mm309at55p
6oF0/8yxEW5CPv6LslAiMPlRG7G0hirq32NBMtuCnSSjor4GvYRXDFPgtCuL/Hz9
8GGUebHHi4R8mXbZQOaOdaL4ZDmjAglu9YIEaKOtDxRpwNck6ZFVC4gIceOpwhlo
dXjsnxBBfhk539UWM7VnI3aECz4UtVJS8ueNa8Eyb/8tGsiYTBXmaiNONneEzJfa
F4XYDOBe7vKiDYfoR3qTDDa1Cvdg6aFy0PiLUIUfW17JXIIOZ9R+5CM4cVFUs4jz
mw0ooPBzTytzu6OeW8eBL5g/A/YLt0mbs4hRqE9KOrMvXeQiTmT63cXq/cs+lpe6
fs5+SDnwGGF1pNVQL7bgxYrcwkv4V7yImb7JU559r1s8WwnQ53wv/RceEDj6p+YG
/22mtJaK6B9D7M38U/xUIJKbydOj3Y+W4XjbkI5HizDGRqcrRJWyyBTvV2pdhq4u
WqNkhYSc2tWkomSM7Qhn5jfp9emu902EhZNJX0zMwuYOEwVk0LJ+yfhLiMQZ+ywN
smRsf9iD7FJYOmhSuGYtR3kdonecnQdt+/toMdEL8ePUOIp7Aw4vxPucohF9xSDX
qVm+NWdvUW69NbaH7fNMUwFttrgBF1CCg8YPQu0laBN4zKeVMCHqB3ooClV463t7
RflV5J6dDivn4ZKDW1ed9igj+mOKziLOj8f26LZ2vk6oYAtsbrQSgkFglAksdji0
j5/4oQGj0iXYHVCm1Hqg8on3W6anw6qsWJu7CEjXKOX+2svgcxCSA77AiFmB51zu
WHGEgEtuZ5MUFbDdNMPjkGBe1AZsaBjPRzSyTvecbJC9kBk9Zu6nr60utnBmAg7p
GnP3OV8YikuyeSdpkCwBp+4gFyJ+bpsr+58Ze3TNjf1P3U9p/t09uulj967l0c1J
Zm2ehnCFix9K1loBlZYeXL4XrM7uDJsDAbo0nDArSCuIZTyrAUYCyIdCLQrkkyrf
1HAX1mXfU1D7KvSASssHNyPe5YAuvL/HvyiRLjv9GgGrtY2wU2LmuQpu2PlE9bw1
Vwc8JDDfDlcHDaAMM2iygpiTaFFa3ZI5TxLrAtNoZOuKknIKgNqyl4ZR1rcgO+Kk
pjD1UddYCIjbb/qWaSFGdqf5+qk7OHgVqcz3AGaYFLVVggip/1t9aEqNXBooU8C0
3eRHHyovODONUTEuy+Ui2PRSBrcT7JwsKhP+qFHCHDMvf9j5+okuYhabfRe2MjL0
fd0Gchfi+IFi3r0fmno6WZfcKCI562LTuhnwAahpdLt5en0JzwndopoMY/2ogfyU
EdZLZSV5S9xNgg7FwAMbfFHQBwAUIwCoXunvvDZ7Yb2+WuXl6jk29gHx4up4SZKi
oeDWXdBa9vgN4G6K5riJN5QrpLG1M17vwiSpEKcyUx2SRqLlngGKueTLIH+tageU
6WKQJ8zSgEaJVrCa4E0VZK9/D2zb6GjGLVns+JrsFfW4XAoZNANsNjplG9VGgDhL
GEy5gPGCUB7jdj08DnU4d3fdo85UfJQHr+hsJgbffBUfT/Ly/zsRZdcZ8zePBg6j
M9Hd07mNiko1/d0WHpcnv3o+ow0srDAxGCysPcsC30jVlvadK9VUrF1ybwqR6Cys
ZRRUSVpnAArNobV25V+E1NqKJZV4YrPBQ3SUYtF+m+PV8SAUNGxKyLnI4K8jwzm7
dQoX+0ejWO5UeJLk6tqnHiuVfIFWMnzvVcClel/48aNkjeJxZ02548d18NJYO8TL
WpfG9p0sAk3kcT6/K0+FqOhe6DDRy4YPi38sYsiUvscd3KsAJSQ2dkygmQ0bTB3l
ZeCJHHMlPUmy77WG4KHatc6Vh9zL5j0Wy0ZJZefkqNfCDdSIwm1fiyauIvoAJcmo
N0eq0C6h8PO4tPVzIBHWigxg45vuN4zsnQ7E3q9TFz3TKLO7zOg0mwwl8/ugfhiu
5J54iWHbVb46AcLHJrEFvSqkMFEwJkYdjD78KL+Mhc8jDBYiVuJozQmLajPF3Fdh
wF8C8urw8OJnx16N6SAadIhTFmva/r0+7Sx94utDA+8+yFhU76nFlmrxHZag5Eog
JpuDcm2qm8srZQP+ny1nwQdqCqLoFAdCJT6WFwJK9s6EfKqVTZAcvDBjbc5c/74S
AXz9kPBXWzNeFfz0Atp0ZprCpfjxy5fMrXYH5mBgfSc=
`protect END_PROTECTED
