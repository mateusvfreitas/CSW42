`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ywVAVr2MvAX7XP5mpbhWThoFsqTHqLsxDns9S3FhWf5nJ4LMMsz8WNCr+11AydOI
/DU3hlTe0Zzqqm9St2tMep4Vgjh9nIDVjjhoHdk22TBlBH8BqgaSni8uevNL7eZX
y5nG2YCEB8hhNRhvTIKSrRbusfbVnVDaHeRTOeFMLzxt9HnTmoHtF+dHH6ZAZCMc
sLrsAwZV3qNNAVq2H9mLLuzQKAoIc31dDmRIFHpi3P4VT5UxDGOzRcDdnqJAg+n3
uZBTmY+aP7vMqw372EQ5CYw/5PEc5mJEsMq5T0wRl1QxM6warbHTh0Hznd+lcJuO
Zz5gaK6+jCH+VdRqJTpNJcJAjZHSnhOCQddAOMP9ISZeySDFbuiDriq+9EEIj4N5
xO6rlRbyBEBae0typVyky24W3ikMSlbIle5SV0FJukldhM6cowH4iDIUKik9xGcW
m/QAioYH/5RPTdkORSKRg1gfBI0J5Dv/WJbT1Z0/lQ/Sel/fVEm/xYQ485AE0tyx
v6kA6vEe5bdkofvb9rZ9UrTOUHbU+FVI5JaGc+YW7zarqnUSgeMar4250tC6Lire
k/iCBKcRbjWw55dGRyssdbiCqGSiWrrU5R078mC1e99pGlqJGH/1oscJiIHb4mH8
OJ/KpkOV7+IyovwiL6znElpuH+lcE2Om7oxFkKIvhyRG7d8eW6zIWiVlQ8BDATM0
+i4C35v2o6ugAems8LwlmuMCmDbrE4Q8Sscnky6dnKE=
`protect END_PROTECTED
