`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
8YWziMcoI+t+BJoI2YvpIqcfBLg/cVGCEjWAkiY93mnupdr/9pwxoo7npQE/t9RJ
xBFyy6O8Y+shkT0blZNzyJ4iQvRSjNvL5KvrfGvxZ4FlwTpM9iwNLwP2Rm2Fl24C
jSh00X6THV9AANe9mlYlBQKelu+59H91wiAD3gswGT+cVbPQNb9z751Lq6QwjH5+
WRzBvGfdzCHP0WoGxtrRfxgzo8hB1kVFbaM7Ms+IMu+sRX+bq7LbQ30cj+0mxydr
+AbOetA4WlbZ1kBYxeRWp7hKozIoo4F5ZbDrrBAoS2Lx6KtrPRJ26o6eoFEqc75l
wt3qGCdlUGcW1OdSV2Xz0sAckXjRhH4D81uOrQXpWXvT8sElDn6ZLaoi3CcBOh1/
aHdyKxcMdEn/4wWmNfMgYvmeNKWYb+IW4ra8rJmz6RkaTTilSS4Sv8D0ZEim10o1
vBF5F/PLjc3Kc66ipHDuOglL7KfXeNgwWPChq8k2eLo7Q0wiyphDc3Oys4DQHK2K
ybxfSRojmfoeM+otKX5WdaWt30HUk9lxRXDR5FM/WIBmxRcAE0TSQBDAUEc4apFi
YtTatyjMqwCrSpeMr0hgMQKp5sbQOvPKC5Xsy6cWYnL4KDO+/6Jwdo3Bvl8AMeV9
HnTQu+jwnoZGDMru5EBB38NTilxVtszl0pLlfi6JlHEW0fW7LjF/u4YxMBYSX1z2
DKbuTl8HyB8z8gEH+kMKZL8cKNed29TJtU6PyYL1Mw1fcabg5cAOOJpWJaK7bLqS
gBA2LzRixczM4AbDfbTWOFzApvedIo86joWvXcBE4i8+JWWwqfc8gqSyqHFEoxNQ
5e1xrwBqW27hjLxDlM89RsT0O2sMxbAQAkrNmE3ZCM5RX+n332jffFfkjr7Ntatk
TssBXeOnEAxuBMzysBvBOBPyvm9CQVi/W5oQ2ZlYO2+FXbc8Gr+zg2gXBfnVFSOp
1OR/B1WO0W3WS/HVwkdPBwg37qDnNAD8KebIxPE6O5aforIxF5Dx1rOziBf68Q0z
ZZjATGMjQig4jZOHkYx/vEti7X0X4Vws6H+O7rHYmrZF9fI2mFDTBFi8VVLTUZJX
opHASuHEryhZqgqj6U14YqInpn/twfBS0q8/5KDEUgtYEDemGwifPncVTQ+ZHqRf
T9TY9uC3t7XK9mm082LFmXEjwx8pCzF5RnisvT5g6/2VIbU11N7+MQDeddt7RczC
RdZZct56SUcsEmOUjSBRyXKLDvJ/uZYKEQIgA5WUIwbPFkuNq7Ci9bX04FfAwoci
IykfOKBuiNhzjTWk4ZuOMLmfFprQp7zfUH9JmjsFxgXRliAO1G3bd7gxgvYqMuzf
JId8aZ8roEzGKe2k10rV6wE9/EGy02NNNuMoUboIrmti1gaeyBcgyLSZiYrYaU4I
sAVF8RV9omrIpLkY2cHnpBprkJPYiu+mACLt2tBOvtswV/bu4yR4g+lwbZLGhhvq
+PnpHmSdnZfx/GxbjYWpAqeJu2j79zRz1NGXU4qn6JrLJHAPRRs3NcQe+E+cWDJP
gT3NEk+3rY6rPGXzUpCooSfPs1rzN2n9oFh1dhJGzOFknLMAxuD9MP3xK5oDVoVR
7Y7tk+N5M5MNS1umWBMmFepQmPoe3sj0dPo9+leJ04AMCVN741U/Gi/YqRTebGvF
Eds+8ZcqwgMfR7tl9yGBxE0AapnvEPJwQv0L7B8gen1SBtdtnPP/PMkj3ENBVicW
/mhp3pbKbY/NQwKR+bNxnIRQx7jkclMkj/BPecUgtPUXK+Hw+mJg+SScbIp5vIkT
6AidkG3USD1njkDL0X9RiZfpPWO14DvZ/kR/kGWYxSQtmBBWqV1P3PHxB8NVf6cF
i2tQuFU/PagRXkZgSvf2DQBZSGmE5jb3QrM5pZF5jkwXmyLk8DxvAf5SE0TuOPJv
4VXkXMsV0O9z+kTAfFjCYpXC+QhkD04rGz/9s+Pl7qPPaEvST9Av7ygdXEFgRF2A
P5fg7om9bdQNh2wy6sPUWA==
`protect END_PROTECTED
