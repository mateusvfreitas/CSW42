`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
iiI3wTHapzr8p0pD66elsXXpHrROuw9QokV9pRUqMOoEV48EVqZ4+2z3OPtZMyKa
VsaPQ2GG6BZEWDZI8P7sMY8mmbi0GHM/zBEEyLYYMScTOfrYPwsjef8F48/EdLUj
cwR9CH04MntUW6ww1/onh4C4P00tLOSAcPiF0xXleeGC1du9JNpQgnxx7bJ2gNY1
PUZKcFfQeu/Hvs9M8+IIEcwi/hhYXoTmIYYzAaA/gJ1MOZbDfSQzqP1Fg0zA5ZgV
snbBjQZHz7kBK52Z4uV9eAtd3Igi4kf56etLB8i/gINm31w2m7hVe1PnGbYicmve
Q9l09PbNO8PJ222TCn1rWL9X8bKsfXwda1xYnMF7n7gQ9rX+AAeOVH0XxFCLZMrP
kSQOQLR4siYT0dkq4rIJ2QW0MHIivOjPntdFDgKpzb1Cis+audTegQl1KU/PtwAr
mL7aop/0BpvSflYrbck8estCi7P31zZ7GPIyeKmuJnwxeR7bKdwlPxBeQM+MRO8a
d8eXPs66e0jR3L3/+5f4aHd/Erxd6qGeDZdYayBxFzvgROjL9NOdsgbfEM7fJ1MZ
EAYjI31PzucAUP0BlZ9fFyNeP0BllqvPDt7i3bBrC77BOAgOmZphMn4yaQ1Efk6m
5OhKCH+5ApLsGrC5pFWJJyr/uovuLnG6uI8NCHAmD0+s4CSJf7BuPaY7yuNa9NWI
HpRmh5odSXTCLwciyI7mjAQDk+PyDj0K8Mv85VhgcWV3ZEjjdCb/SVpHYzTFcauV
2w/uqXyqk7sipIy+ILET0x8kmunlb56d2HheFpH/IJM6/THoUvED7TWkvhQkJ9m+
0695+9T+ls9hWqGv1JDM0GLBcrEIn+8WMxVJToMAlu2s4DdhXB0w+CxrsdgjrOa/
iG7NlHzNE/CX2XcaGdFb2Xytp6ZwT7tCqBbMsiuTh5kON9obP3GF9cDGIsrphPHH
4mX+L2t4ndOCWNDtJWkmj0RjJs3qyQHkQbRDjMhYj4ysTCj7YEfXUD5uTmj58EF+
XQR5qsZAvIaHdygLcespKF9caMZIQm5yGT8xrZj8I/v1dh26897X8ISmmqqayPkh
VPp/HskIvLPZQRPw2GMUnaBHBvhG6G9/dqGS7Qs9Id+8Pe2vEEVacplGKvDgLfLn
cQDNqjuzV95CDbznW8499RI0IgP8jr2kj7LNlLmm5RZh1dVSpAlf8FxHh+2d2baG
5omJ8vR0VOJQq7vorWPMIRkgi/p7mpPETILqfNxGWGd9ybQK/3EAuZ9OcrfLtAiX
g0RASGVs2uWIdqqTDyz3/7vn5/TVFZ1DgpsUdbYuyr1iCaPMw6k9YwvnCftj1iiP
J+mXZZGzrAVEvcDm/wfxng5MIsMVbxTdJISeOdlWwgx7hRidZtAwrpJWPBeOwuR3
wIhNbVpIRCXpR1gAo/r0o0+xCqncVb4bzlWFfzu7FSbibrufODPWiU9q/V18Zqqh
hQYbZGMWjHQ9QnvrkW1l4Wb4IjJA2oS4pAedgxkXiOnZ4DRbQDXYyQ4+cKGYAsHV
uLNMoek23x7inLSRBhgWTnDTksbyPrFK+S81wtRs9xxtu+9/9RKV5SzigrD4amUW
jF8Z2MtPrTgvvixuWI6+oUS2RKTQ6hYrXcCDmAQE+9eQVshxpU3+atVKs7Ggns+k
d/XuUMqnyUw3vLA7oaTY8wGJbK03PDGDahbWZv0N3tOrYB/VpdEpxym9w38NErxR
RLvqcr1sgdWZreDt7u2BzT5l1f3xKGhuxz2koP7YTdoBqDtYmmGknQWwS/dyJdWK
JKlo40IDFdHs4iyb3W1ghdczpqCXd9nq7NR0VJz5EJ9Z4GucPuUi8CTU4vqQnID3
n7uAGK60TlobTFoCk1XS41JfZkVNcrsYVVIlDbCjBJXtQAowMzQo/yMeQNysrMl/
f2PEhrA7zsL/La94Tm5TyLolMSyByzEauVO4i+IlozHjVttgRRCeXgCdWbbDcJW/
wu+2SdlqlB9ISAU3TX8XOOV6CR766aO/6B02bEkevpWcgdeD77VcPCy5O1nJsfx5
`protect END_PROTECTED
