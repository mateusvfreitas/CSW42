`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4qNGwai502ciDhR0Q21ClIaDFNC23vbMKKYizq+zWlcF33B3EGWyUaatsHu3YiqR
zrtrsCmSyG3qLXlQ014qwx+iPNe1sAMSeLbeUGPRYQHf7ydfJZpE5nBUQHNph8ye
fRz+p3GlUeJYllNUH/lmrLVQaK6WNmckVDik6TV/T0+lF188qwXZMqZdHbOjmWHZ
lTcBCf2u+TEzUO8BdZoiAuqsRwum8hDiR1jkb4gt7yCyeS9SHWzNa9Zxswx/6q9r
X2HVVDWE8xnmhwM9RJ36pGdjkL3vsOp8aJatoyNsFviS4LyI/lAeKV9loPsmdatk
AsD6/oI81u0j1o1I7m1pWH8PCLOWDYYiIkLRaHBE1GqGf57QJleZTmdSC4ddH91s
34ttdgQWkbpILGx21oWLK41ZiYAgvqlWZggbQNGQNHZRBpPmPUKWJPrqbMEIdjea
yok/Z+n1Fx6Ip5QKI398GlMI2/pVUDyrqyUks1m+2sOpxve4A19YYXPwHWTLIyab
kZzIfcYSONu48R3OZNBVLvNnq4tagqWjjSVCJecRXw0RdjivcqUHgA9rpETyxVAE
BppNzNCdP4sstGA5iVBUreT7cJCpi8kUB+ytZBiMLQ53Cgq/YAs/H2n6bp4z7Vq3
y6Hgq2TacWI9vlmy42pkWhEdPoWyugRKW6aLmxR68+/Sb9a6PXqsvj9s9BV7Tis1
I0jPoUcTlMRopEx/dTNidjdi24Pcr0me+8XZdHIU6eA=
`protect END_PROTECTED
