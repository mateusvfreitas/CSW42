`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fcNP09NzybpyyvgVDTTw14tyJyA/k2kmehMmuMRlUWFaH1scJdM1m/ZCldMRJCs4
K+tM0KmwV86VaGlmvodd9hz4vSYjXUZ2UBcqaOidNQP+Mufrd112eFsfpO1yJnG3
wZ5SPkj6Co725m/cTJLg6QouC5gcVaOTao4zBL5iBGep+HGW1+evBrUNiHdxrZiB
JzxBiJo3gsgxHMLDZPPxvooPsBhtipgM0dls3rh2NWdYg7koae3pDihzevnDDAH7
zL9jaqQP4j+sKAKixAXh0DaDqmFey/QZBZSwJxVKpaFP/C0XuxcTk2aBGnTszkjl
arp67bmwEv2pJMKgtEFF1JDl5BkKdEB/DDHDFPJG7GKcRaKw4qMYRr0FcIQ5ftjp
I2An56EpbGtzS+jEvTS40L5paUcyvsFzn8x2ZHlrgnsIm1yaVh9GpoYE+pZ2BXAk
KLRAQXzwVklAWxZw339WKTOkQiyJUANAJtesWyZeGb2kTMdg9tBZe2vBKEjp1EAl
uDw8gJ79MyURNTlQ39fevpxsuGEgHol6MksUCfqxT+wCQJWIAX6BISO71JHXl+wD
Cieye+2spuV+GkHVMCXDX3UaylX6qNogo+yH3US0BCCx8e8B+wrKxkmLKQEvNNtk
3d0UkykIpf/+lultT0KtCOdtxYAmwTJhhCwEyrOkPk6szPvjHlALQdd58MRq5yMy
rknZ5IkiUCvLMFKNfa1gP5G/TCgMzzbIbc20mvy6GddYjDeV03rybz8Qsrc3cDMb
Jm+6ZhazTtYg9FsDVHtB9u3kiug16weBoxcwH9oXIuoicHlH/ebRtRiwJv0UxFw7
9E0A20KZpySUcAPN0EdxBWJBVPa3oTRLedyPhHFwsglEO5rOiuvWnwIooEp5oxpY
K6yiX1XDDBtst7LOS3hdkBwgL2ZkFJ2rPIztdV0lbojJe67BUVBrXHAe6kVhQKoO
1Iq03Wx0CrRrDv/59BrLXLxHQMRFnJ0/cHcbswlCPH3HDqyEKK4JMPb8WsBpHFYp
/sFV3n/0GZVIfxUaSDsoIQ2QA84j0vy41vzrF+LQdPrI0X8l4CuHW8vXj19LCM2n
dkNLDxUIiVLnQvXGj5RAOCORbH/9BiOxjIgqs8Q/JpBpmAw2Qa0+6FcDLtEsoqLI
4DQLziWG7kYc6v+w8rJv49iSNKQ5cgzcAeSeULukEMDHxpi0VQ/l7WbMUi2KzAia
ISOOPZtLluKNReygGSjLMpNIyBsnoWpZJ1NRd9hLWYM0Y0bImZDKR4jtvnK55r1d
UNjuGJ0tMbbr4Kq8tSJcIiv5FmQxQddPvgIBZQC0LxEsBBqZXLweWcdzTN7rt7HQ
rgF4Iz4qfW8fr80SZaeWh3Qxyv3IU+of5WZ3emUQQKRXyAvbRdFoNp6OyP/T6lXk
RlYL5ReSuexgRqm8plUT/7kz0vtq4U3g2KBYEx5ep37ukidxl0C6DYfjh6A7kVyp
qG3BT1/xxxAam3/EbAy+4Sc0eYrHH347jAXSnDDsbGaewTnoin7PeGM9HzlgR8k5
6pWv4ON9q+fA2x3yLJ8rwFQkr9nklFmnhZUguvpMDmW3osnsrstF7EEua4lh0oC6
+IoJ54LJskVbng6AHiOYN1C/0zHeCLNCSmtjDr3GQ6McUEjrZBDXkss630PWOWmX
MMAyaj760LrBUvyNJAOR1msJMboGyLrn78aoA+sY8/MeE9K6gEjMDhYKfN8uvG9g
2mc52UviUwULdicRfR9G7+Kgd/Gdbjd44HBCWTbmgmLd9nR9M5YtejJCpQmQi9lp
EIl8NIUaAFhaAkOIaFVCXFKR5nPi90k+8Za0Howx37pwUsCQauRHCdSONvSuwEoB
0gqkxySg+vutxn+K8CMjXwOg3QK/RkYLqVI/3m1N7SjRNqi087o6BDxfxMLcOJDt
N74LvjFr5GqapqErx75nf3bFecKKfByf+iYmpRMcf2jTrJ5dYI5CIJSkMqiV9hXl
RZnWVI9hNTBhhj+uvzgHlyzX0LnmCzIy8QilwLnNsXm8Db7rfIHcpd8/ZWZdusRt
Gie7/bVcvJwBKCh24HpQ/BVEQ/Ku6yyklJgA/ZsbbimstLA274Rmbf5zg/V4Vp0y
bcH3rs3don16GsmmzgOLbJB1dCJeNxdB/050RFdEtDDF2gvrraSbF6m21PNngq8M
V+jnv9DB1dTPHWh4LAc0RftFX/jduMlzqNZhBjMRsCnPKQRrQ/1ueMGC1/EsYuOJ
P2Mk7m9csSrWGUzWaD9nuZ2MYXdgdxbEHl27ABb5DdylHroN27QaOX+9OGV8F5Cb
QsgSzoMBrmWhRRif8y9e2gqoMoad1g9YP80PQ2IqC2EydlpyVSkeTYsRVAB4wGdg
/v7NlY0zddZfTm2DyNzXgpTfna/zd2LfuXWU1WHD4U0cLen4mukjEsNqGn9ohQN/
EYbKbzbb+Bhmdoczo8LOTSJvtPw8CLH2iDK6tosJ+eMa9+2ZT3ifdkTgRghxt3X6
9SpaNedvG/4AUJyQruDq/pUE8EnBfyfaM5QUQxTUtHxpVQykaeogjmyimXvZkoWs
5ZYtMiWfhErPMV4VwR9hi0if7a9VJ2figmVIF+z7mlcgvY3TCuGkCitceXOLdsdr
k5Maa8vh1PGKVSVyvJqdgk1glvuo7Qnh6qBc/eRosZyzIdZKW2S3aeqkr+ULC6c+
93XIHQVYJzFmx17CCrGz0eC+OWyPSFs3ZGngfyRF0LHiz1zKs7nYmZceU0bU53tA
SF12Q+HyZP2frxqJDPQ8vRDmqUTQmrBh5KdPxsm0kb3EcKENdWGwIgvMD4dT9Dv4
HpHKB5emChnRepLQTtWuj9kRn0LmAFzHwu+F7eCqjy4uFc6jWeaKtg0IS6xYOWr6
SIhxwzMklaYhogHAPFie1nj4yGgNyDLTUeio7w7sgP7KS0Agq3LbtSznEyTseiDD
gYnuNp6vPIQti35oYTu6/CE3U6p3riYAQxXaGNA5ETyd6o0SpkOhSwJqJlgareeA
mCOZlOIaGMju9Jr3SiH2AKyzioDoZj6k8kSR06i76SMuRsi5U/CCRFeKVnhUM6gp
MS7UgwdnYYP46U8jbliczj+NWyht7DjA1u5anta0unuiz9dEnlnvAXBQCJvnyW/Z
JBJkvHbfH6D9SzG38kY3r2f4LHYABNdvP+DedoTC5yUIGr5/YgMvjRBs94lvYFkh
9RoGo/QZk7b+H8g2ILR8FSwbaVzYrnm+navrCe6r94wD/r5Vl1vOXZURte1hopBa
7BPLb0YpatfZxocipYVJBnKS8ClCLqbBVn8pFwHIg4sVS/PJT2R1Ghnfo26x6/4/
TFblqz0VjnmtbXf/bhvjO8EJWZmQYPmtDZoe6baxkTJT+79ycKhcqOHN2gqwQMqK
KFpeGoD6PvzPFP+YEXkhMwCW3P37vqM1Wjmb9yFZoXGLTfbuaU+1GdTngW7v4l9a
wgwORxc5Ue9DcXg8vGkXC/mjZh9HnwAnIIDfe2GB9xAMQ9m2u11JnmxXsr2B27e3
NLfPfHBgxm95YBhPWTURL7OMo4b6XRgfbr0SpQ7BrwqAIK90gCTGWoCmxapCZO1V
Pc6Sbeulpzbz1Lz53O5WjACWmeTt+O6VgJQ/XqxhQhuzkGxaySYSSlBcGOgs5fRX
B9/fncpD4j0M6SPULkyZoScyqZfvsKIMSV4LNAtFMOeRSP1RYxY+Ou25WX14YC0R
Op5+/6ElUrIBhdrEaSQMs8Q/g/XstATFN0TDH1AfQudhJhXHHF/mYRu1rg5yC0h+
Ad3kZdTArW/hmbxPDSiP7BasK8kNCfV37csTm+p4Hx7MqglRtDsb1kSRMOqvGn9o
WHCH7QYCmFDsULWaGaNXoJbsC91MWPHZMhPtcDUjfHuUkvkdhFBD/8IRDt/cwpy1
Kvap4CvUYQIaZldwoXtg6ug/OzRS6r5dBUHQAS+JZiN9nOfz9zLOzjjvCE2D834o
pEaZ/p3fCZOep/yS8YFPf1Mbx0B1sWycJAj0UngHBjP+wexEGZxJdjHbEEa5WiAY
8aZAGOoWuC0VKfs9+JZFdXPGJR4dSe5TM4iqc8IEDyy6HEjzwENLfxMqZPZU2n3a
sgV49clzlmGhUObSm41wZhwi60dRVYYb4gV2a7tFK5JhJ5o1In+/nAS2pFdvmT9Y
zuGRr3vS6CrgyQ2b4z7BBtre60g4M8rN2lBMYJXo3PY43SQcN3ppEpaoBQODVf1e
MUanfQHd4GpyLHvlTtWLpU7qfxK08dHtxg/6sIERnrT7OHSoRHLZzma9hLSPSffG
/bwze+CGsidZ/RUeKzSiEiPQ3whG0l13GyjwGON/OmPRLgZVVrEYtnuIoOKB7WdX
6Ge9FeWPLBtWN5wt97LFlele9ojim5H6bnKhuGriScwXLrivs6xXrY2Tcj0rlWkT
yZ3aAP6BD9T7qLtuwUfri7TkDzylHfRcHM9HkXXyAQ7DIKbz5xdDNAzXjr1i7bzV
02KNkItk5M+vMazLXyL0rjP5IxvqJLjsbm7R+eCUhW4DRaUTY23MbxlGihexgVLS
kQ9qOJIFeKygThlN6Tp80yfqGF1OUgtUHCcCMLoMnC0D+xvTwqH1foFRUnmCDc59
UCBuSBBxWH9ekA3BJYvpK/eKiL1mfxRV6CfoVIpE/xp8UDgou53J357mtYsY7Jf3
FcGoKUfMOBBcU6xZjwBHmcJQR+jgYsNf6hdQa76J39eJWVo6fCBm6cIabCIQJ07f
e6+KHseYNBaggjmO8ntEelkKf6JozD4jbaUCopbln9SEhCxOwRD1ii4FE/SG0y1N
Y0g5nI761RSKVseqnNK+r226ozLgZ27o/6hx4qihFOmH/8Hw+dsptTx6YtxOJmjP
qyiChCGZz+hOQhZgGJgteYE6bb7tX7nVuEQslEh/tMJJcsmtAlfH8PN66oQvFH9h
ZQAYmBCa87RApU0oSKWmmt/yc0gPjZlu0LcekDE7nWJYgUooU3P/VkxGaEXiJaCs
l2vR80fL2u8kasGaCAfwUCZVJgPDIozEZMrjR27D1DSfNLXfBqDk0QeGYY0mv9Xk
2AhBEtiPcbFgvLw8+4ukxGaQExTZgBvUFUl+bCaFzN2vFrZQQK65yv6NqOZ9aUW3
mUnn0LNkBZvFnMuirnynIiQyrtS+OY2Fz0zlVPg5vvR5GsLjfyYFzw3dIPXtg4dU
zuh/xOrcoUNVyf+NaWljjvDtK89XanpSy+Ch3Hd5rotqI5DvxWufmwnWy6ROWSHS
YieMwb9oZRCrzVM6jvJB+63pf+nIFxN+LUr5RH8LCtPFd1bcBuWNKQtZrvGGcutI
ON9XzxDOOb95v+Et5jwjSMdBdyZpqjl7cf7A3+j0jVFBnDyIzfhHEgllRchgzqab
Vdoyw6aPD7sDY1BM+iNImUMsLLc6rvSKvbNcvW8JVbbhX96q0wt4cGtZZHOkLnVB
Tw5/uYJdgdR46BpzCnXqD1ioTfEkla2Mx72m9UpvGnRqof4pQeCaY7VNlUvq8o/i
kv0vcMT1D5prUR6R83GIWJx4unOVbuThSzuWFnLrQvTyeTc3V9GsUj/TLWptbevi
v5slCSf8hg9AH2TRf3vqBCoXb6iBD4bv+vr6KrnFqTHWv4tmgLojWCd7TDUEMDvr
pneVjNDBC8MR/+3kcoLHmJ3NBQYaU/MIkfhKR5odkrzrair2+/WtNCyYxzGqfk73
Vl8hdNUwX62hM4qOYKzJCbwytM9HXgqm3nKN3+u7KTlSdfj7PoiXU17OT1ZRLS9A
eDW8/zPAp0KQR8pJ9krXoaD3SRfWoRiDW2bcsG6ZxVdejLA7/il5uoYDhB3wamEq
FhdNODM9Ah94QDkyiSp8+3eJLRyir86q9mj0JXjFUFYXC96O61aHLk119EwAO7AI
ohGmttHgl2m8Ed0rLdpIVFNt63nw2VzJ2iQiv3+GkkVscy+nu7UQLXUI67Pn9LsU
DH4Q8JEQ0OovtigntVUR6ubBUO0vlyuGn6TaWlp1Ec/zrpKO2kAW9/EKllq22P4n
xnowJfb3c6jhVTan1CyMONFJC4Omwed4VH6/PZZwRTRvK8EVvRz4THch87pA7RI2
iPvHYSpeFZh6WQdO7fbuWbggymbHDCgAYV4h6d5UlNJoKSwt7++JH+PlQ43EoMFj
wpthj21PIqcSGU1rfvCU1cJ1B9pghZ50iQqZw9gDcZjk5Da/FwpTIjOIao0jbP2B
U4zhnNRyfeGcrtIVq5Yj+OfQYr9NxUvnW9JwxbBkj1f4MWJe3UBrJUgMfRqNLDtG
4mSo2AHJ4u+lYt0uMamwjojSUZtyoogoLwVGqX1HwtC+P/E1gb+gGlcaPBxMK6/K
rIrq461zNrGOMbQYiOUk0CYV4qyWc9kb5E0q5qqwZSBC7PyxPPINHKArHo7wblpg
cycm9AsmfVwXGVtxEVAJnDSbbQDyNxr9bSuxwLhxsiNe0MiToo2QMwtSKsBcvkmw
A2g/ZCIh2E/XzDgo57vjJcNP6Lzx+ojJnUQwzC2rTo1+jNOn5FYMUzaaUfRIhleR
o8Oiqebct1g+wmI8e5xPHV5XBlehCs5cpQDfyxeL/rJaDE1R0tPSFYkr/5wrhn4T
kvUAo6A1fS07UAg8oQjIqAUm1OQRUbE/inMPYdAVW5fwDhqxXU1/TM+yLcYqDp7l
NYiySbKdnvehi1SobIkgYMDQqhBW4Nrb0Je2610nKiGfLI7Rbbe3NK5hhkTi6RQX
4YGefJcsFCnod+NxqVxjTS55cr9md7dI4IlrD+RhTlnq6mg3QAjyBnceoK9SvWPe
88PKClO6GvBFNMcHSybaxZ37NRmWWtDcAF5lfjAMAoW+bxRn7T90KJisFc4wwk/T
5aQ94u2WzyHSAk6ABMRzY9bfI6hPuGvKDNfmYZw66LR4QdUD40FEVggNNSYdrzvj
5E21bYZNDbjo8myp2oOVrSyH+Tq+jahnwuLS9Crwn8z610WaNB7Dt4vdrPWnqUQu
pcj3N454iNplvYMoPNM2IjlnQHbyzIkLvVyskhqhHRiK22B17tjmvVQGwj1xuEbm
wv/8FEpRrnhikgIzRiXmsfl23VsiMBfq7bspCoBTUhYYllr+M/NIDErP4enrISEL
vYujxl0c/Dir8KWOmkeZP1YtXUq8+0aMTBRdXx5FzCj2Oatlwz6B+IxAXPNLfTwm
luLfkBTr0LGnSCbjoBj+6fpMEAoJRA3AQ/gD1qrml3x1FrnkcZ4NePuTI7oDNxC4
k67nb7f8Ywn18mV5lqi3huNQCXE1CBwB/T1rAG86yfeD3QrnRn255iZR8WpItOeP
xFPvfYFqQ4Vh2sNF6go0SSaUdE1cV0TvgYrAGkIHJCqDpwWsvg6Zy/IjJlg9elvd
fbH+SVVulxeX3uQ4OktnHhL/umhKf9ElCNJyGE2uTABOx6vOwNo4SHM+KL99wYbJ
BsScxRua93CUc3l271rxEqFpIa0NdSEiWnA1DG8QGSsIGAhpTJKWaVklh7G6QmfJ
S6sOFU8xloexRZdNLiVx7ad5+Kwe7YFrwmwkOMQU9O5UK8aonGkIX7CY77NKDLNz
vdGpGeXduu1jIm9xIAL4lRSLzJW/8ijcBrlYy8Wvk6vI+U03EHSEdyrVBY3+yP1F
auqlC0u+rNHZ+QORYv2hxt7gWk7PGD8/kE29vXR8dqYLgSWjsTeN1ivtUoOCn6Zn
`protect END_PROTECTED
