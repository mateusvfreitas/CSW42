`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eLMJUe5wX1Q9quXUWlZV3DVqppBF1t4P5ES7c7oXe+EwTl67FhgAUcWTlu+jm0Gb
8qXJau2DH2SOOZHqr1kaV76DZIjK6XBGZqBMHYFz48hHSj1FCYkWA6BlmvppcUd8
lIEVh5qkLMQYUDUxVnDns5XLCs/K9g4n0cLC9x/FbeYQgogkst461PBq/2JVSRL8
hc6RZyiV5OfGGNKULnUcOQJVUxxrqj71qVolYXFbefnpQW8XYLewNKwSPkOfxtB3
p9VxZhbojOtc6ZartwOQfq0KczHc1qSdUysWX21YLx5hIGqUlOK3vUZNkQCK8lV8
JSpgQT2Yb0InnVVUlMImqOWOWYJVO1q1MDnY8J2t0NwuENf9bOtodkGgMgEFjQvC
MMtNhkGfLZ+TShSubmDKijMOJjeoWCmI4uSuy6kx29ksJdLwATHbOp1HHnRYufVB
KKijOHEzP7VB+iAJAoEhVpkZ3MT1XG+9pC2t7OrsBvKSpObhR9JhZaYvhaDR4UyF
xrXcWEhz58lYNVcpWvtDe42ognxXy4Ib7RFWZ3Fl1GBQHC1NKDt0U0WIJqgB+RrD
X1LTuGEMrooAqAJHgrtWM1zRwOeSELcO4qmhCniRzDY+diJOsOi6Px4ZMz2+aqYj
VARl0h+tsWvYz2IU4T5W8LYph2p5qS/SEKOEX1ZnolWXLIhw6mqBItgdysHqHEs7
Su8Nj88WyLtP8JqwyrHCK8yX86uJdJ6jYKcIOQT9aYrR0wLwXYBzQ8GhTsjgL4Zw
+s08HLTpO+7TW+YwibL0eFUgLJsIg/yXmgQQsHWZZY+gUwjeDBhQtgIle8w1yIWh
g5+zmNG8RRXDdG2SkofD5q02/plBLY99c1DgRF7hyo+Wm7VC0fDLDJkT9X7ZnEcs
P9HdjuXAB8zyLakxQHdjrI1te243+Czy1wwrnZ4Z6DFjiO2gEahG8kO0DDlOGUQP
nEXDHOE1aPFE75+FBNfZB2GEtslHXM/NX3eNRsuleFsy2BLnhHrxpyxU3mkIs2+S
Pob9w8oGygqSaH5nEuctZey/7NTE+cNPz5BOMf4V4R86Og6jLNvj0tnnJoHM32R8
9KwqNC1KNed5FslrxbQ1ankw5bPea9ncb6fTxifZclFA4i9xv75qLesNXDaTzzVe
diNybM/hRaoDZWFU49jgZatw+lo3aAPpIyGytBK+xMnDWPkMJ59ffrwYaxm7JIFS
M1L1ml0DCDr2FpuJY+xRcdNFyzwYQI/Wbq0+2Eu1K9BnNX5Qr5mL0zQA5eXz01O1
oUH+Xz1NgQgDfWI9bi3Dwya5saixYt7mSzSbPgkjja/Qw9O+bytbstTb+/VUU+Bm
SDhsvUbV2e4jWV5N9abOdLlGveeNmqB0XmycCu0gpoh0u6F5owoqQy8sxlDM2PWP
z0KGRr67r5Crnivk69hwTWw7PV1AaN/j0Atl2SeF7bhuqWZJYVf1bFslPzBoR9Wd
TOHcOKlmtOU2tVjzF352RS6nWye6PFgIE8H2DDCN92GviH7pBnS9eyS1+CR3ZoUS
7ZnmtlPAQ14KgMbcTnajQBPGboKDXKsQdFN7cwYnIYJr2Rk9R0F+YSH8rUf7FAdj
U1txbd4LuzJ1fSIZZmWXPtIAOicVKouGGe1s2R6rD6IgvLX9QrYLO8NTFYpAuFsH
yU0JpWG6cx6xOudSvCnGphj4m4dL1fFx+qVJyQbKNlO+enMICJUI2ZaeJph3UbNk
aI85AlBjQ4y9FnW286LAEN7fRCCk1ZlDWb25NiOkDnU1c2s693Q9tZWazMLJTdS4
k+pDSos2SxvbZEBRBjqXDvx8sCysbcweT4sESVpSj17UXOvhvxQocjc5XNUZokei
mdFvIrffRM9Exwivofq15knzSb6NS4CKQlpmHJQeNLimJa9i005iGbrzD8o30H2v
O01k4viIvoXu41mRWGuKkoqQFVBvDZZdfSL/ifYW1FgIpkseixe33bpgRAO38fYc
ZCw8g5WmeghkvR1TO24+Kfr0hyF86a9AJKwwTcTUNz9nn4ugfaxlV8ZZZgToNI1L
KUsHCqiDwh0ltbSHo+Dhcs3Aq0rcFlwsEOikdrfa8ktt5ysCFfe2oUD3rwjYg2kP
3AYUnxzdiE9BDU3/BsF5rR41EIayAgr6Lrqp1K2L0VerImwN388BJqTONe3QXqMF
p8IrYaHf+RPpMNkDPnkbdg/6hrfjr48G/GaNj6jDiTJs+x0PhQkCjYDk2Y1NhkY2
vIEB2vFcZVAjdI7RRnb8XqezGpZzxrWdVF9+hg/P0+ER/4rMmuWYSKHz2BZGKKVX
b3lM29jO9iG05TBWdPBMlpsiRN23mhtz2/Ni8kKuI0XA0IgYr2N2Ym8geiyI5y1c
xbzSkfxt3xVMVdEfgUu/tdIGKDi/Qe8VBkAlczzMWIGQ0ETQSMgrVxTZuSfyHQkr
t6V/F/MvH2whP3t48G3mIXbyCSlKTKf+LTO3Kj2+mcntAXWveN6vKFAGC20RiJ55
c4UM6vE0Kd4+MFXW8bEuvFN3tsHKYWUESX6+QjiVWdv1KTDlwPo+6YuSNKmKy59B
Tz1bSvPaRlOdYHzFwtglq46yhJ0jyf4FfrX35cU7USrDHCOpY3xTe0bpp0WkVxaj
yh91jFdhOPPCddO3b+e9OCvGFZEnnZkj89dKIy6ctFsnwJH/DBy0ilZ85zMBSrQr
6cKhScpWpu+0OKRqGpRQN3bu9JsYrIZcuukdzy948Xz+hJQfG2/qXV/6+PUUGfju
V6L7qRMmTinPKj0atrht/4RdZ1tBGSXsgmWxbFkyxi+W7B8z5I6bHoV4ktUpL1GL
bNUrkI+OBgBD1j5VIIiR6Uug8FvXGk5QWXiXxXgUGoq2MREEacqX4tpESi0X6Pq9
GW3s5ldWWHLVnXaVBpNT8L2fCBjV+ZJbXhEGCTUXrVSkePILofzGCaTsMS/bYwcJ
Uzs0ztYvcX7nfhENg3JhhUuH3YMrl0ho/01S25Gm4gs5cJKOVy6IBW5IDdPcDHCH
zrqfW/eK37p5Krs45JPGmQLpMQPtauD3sqeB+wlvT120evVT1L/JNTIgxiB2+5Yg
fetq2fTjJu4TVuNz9N3GhpmekHcOzKH6jlsD/ng4A7UzHLuSBjDMvx6o4RavUo4Z
3cNm2EaI7Qb/XjrXxOrRAodPVwz3PTFYMiuDR6ZA8++zVAqgIdSfyBMozXIcUbz4
S1HWjIA9KuxmzphPqs3GfPPFRcswUUGNQsE6I9KQ6V3i66Qxt2MpcaJK6BpYuPrZ
Q7II+a9OLV7Qy3N0Aq05vIisI2AjWukrXH4x3MnQkHkyChRWBQQVHjtPQNOqgRFG
21quuGo/BTmC1y7Y76kMbRJjC+hUylLjAK/0YNt6U4n8N7JR6L8Hi8N5U3e6xPPI
vov8J0ULGGrkLPZRveqcDouWkW/p/USGBcfv/l7GYBsfiJP4zVsE39l/+IepCfsW
7C21pVvoPiuuUA6Sv7ZgAEAmSJ4qbzB5dEAPE+oOv1NQCW77zRvLPbChoOwseSKz
UPhtXMsNDxfnLSsdCvH2yecK5qHpayUqGsFv3GO4gkh0veuXfDxW/4dafWM8Z7Ua
DrcHDratxsOafzYX7EAAZWIbca3oDlNrJRby0RLkaL9cux+4igh1MXvp7SedeZD8
kUWnIDxR9v76cmzgCfBbt6IBfKJoe+H7YrbQxucdsyAWlqBEJAR+aZ1VjOuJuHRb
fllgWlZnZ4gsjnU0COmku0jKeqV5G011sgAkM4SQ4sICg4DcGQ3wCnAlnLy48Pq7
cIq5nbzF5USb/na63URt5gC/uf0+g600CHQdoSUhdBvM8AyslyAa+LlHeBjtZYWJ
JcYKiZQVxr/rg/0A9g8DvU/mQlh4EQRfHnDBbao2swCQVZ6Mw5YicyL44WPn3UlO
75JQwE+ECztMvXQHfi8LjsYa8N6jyg8ncDLr6fKegORy0gWrYTDVifJgrwa3wMj9
JUZJlu9Zh9i9YfQ4sTkfnNwFQF18SraF9+k4Y96LBdAsj2aQw2KEzBth54fFvnXd
5f6Iq82vRiHYAu2KhMSaz17ewXq8KYgUf9UCwV7X5cYuyW8rd1Ci5OJEo816IRm4
+6GJH6GGv0Wfn2NI3DjiXBIUUMocampi3FMGEnGuWayRnxEpZDm0B2p+RYBU4Keg
dQzexrkBPxrZBZWoLSSPzhEudydkOfik+qq3dOkhQH6mw1EM+tLTr11sa2/axQ6+
srE28eCDvos/jZAWDH3ndPn+5Qyy7Vo5watRgvSB8HFx78ulD2zLKgB2j2W/3qN/
GzDfx5Pk6+XXDlWbZJ0WSaoGrJaQ2K+9s67VGs9Qh06axo6hwsgSPgzygYxz19X0
ilqMLxk9zChNgQoAbjup7k9IzesVBL1g7Pqyc8QGkWT+ktSPkL1r8H1nNqv+vs4U
uedq1bR8TP7O1uYjFCG+yfFfwC8fMaBqheB9AHaN4ASGjA8sAQgWUzNEmm5ti/qg
Jv81sJ8dUCEyI4U1o2IEbyzk5XdC21AJKmfET38bKkO/16ef3fJSItHdWyJcPAQ0
NfkmjgjncMG2pM6JH6RwstMyV1nVw6e6rV5PsecaFzd7tQzTrxv+SYy1EyIptjGG
Ss7nEH5RNeca6V4ekb0UlRTQD1vXx0+RX/MOy+ifgKnQzzBPUYJMQXD+LJm9nxPQ
vtnLXnrzSNfThoO+bl2AEPmlhdq8lWluh0Dto5WOqWMXzF7NuxTOfwYh+/mt0puk
S2gawv9r2X60Jsu+ToT7lSI5ZzMshTlg1x0ED2Ynoa4cUFRBywPeWxHzruIjSbLC
7YB5FwN7vSmlWlu/b/+sdTlj7erBCQGd36gKn6+uz4JWMbjJJZhMmYCdm69Ch1Db
MxQMhJQ/QVv5ZPfMx7+DnGvK2LZ7EgKGYeMOMSxsuybNsTxmI5pK6t6yVMwSxEAg
0IT/v7dDWdm40ZJxCHjgoUN2IUbuNGk/9xjDGXJ3Dz909Qk4mZc1oXQTLrgVks5E
hnieAfnexPJ98HIWaUnx1wMc5a242dMgB0JB9A3/fpT28yMm3Ow5yKNYtzxVNOvx
R+IKqaXZvMMMxXqgy+Z/YjGx46vACtlDmt4Jxf8gE3AWdwaG6BS+tHtvc1JWe5g5
tsjMOS/XeONYkKsgarpKzENkWsOn88tHCtWC2poVvivbJeWvmx2FuG9RCTYWM1DV
P959jl3vxAM6yPm5pv26+iEWv6XlpgzbzH49WLgzI0+PI1uhI5f4+PgfvA0fxcfa
cFsnnJXBhQlbcOBHFdVIQZwaDrnma0J0ZE85hYJ7X3u+2rub4IEAfDCNsJcVrLPJ
SshFv/bh0F7F12G4IzqoV18CYLUh3pHG+gJYHe5mtlcESehki5bNdtqkfTRtic5D
NOP+wWCK9m3v3nz6JV7PSrvWEz6KqL+fZI4g8Ad2kofPadz8IMVn6Knq9FlUNrmD
ynrjhJxiHSSo6zwiabK9eVFuhKDkVjYy5yDx0v9FOImM7kHDP0U/mBeedYZB6raI
megt19aOsDCLlFcVACG+VoX+YWlw7Y0/0b+nS6rRh+KD8d3GVk/0oDqpf98pVswy
SOcTgliOs4btj5J+GE1azceOAEb+JlPFzxrRrICEaacEuIwq74i7ltp91gF8D2Cg
t6l6W9zZw+AKrFcvv8/qyCNi1lQejfU76PcNvKV7SVBDQy90rcNhiReOUsd9EdvI
U4pxo1FFCgGHeJPRr13619BQfR/aBU70HmvMwSxugerW7I5O5xOr3WyZi/LLQCBq
7HPkORw2AgKEXyCUmyhX3wtTSvPRlPdbhbPQCZZhyyyDe+aaYC1FMlk0QWPyESwd
FKl0ucanLEwdTGwAG7x1vd8H8K6CnCNwMsvtgOiusDiM7DNc46qp7kctTdl6vjt5
uD8yugynZ3nci5lGx9KvtCwL5I48AkqDQt81+5xyJC4VoAecanU3evrPZQN3Qxki
AasV8ykrrCJ+YeAkl9L2YC0dR3OpBN1Ltso9p80u6CnmQkbwal4Oxzz4ElE2tnqs
6GD2WLOcZXpnAz3ow6hGmb03606ip3hRtybKyAFCQxoqU5OwshqoQX703fnFkCzt
lL30RZ3qRKsU2XcZRYe1SnRCTE4FtJEXlxGKJCRDLlWg4dM4CeXNFPj3SSOB+ldw
Q6cOHwvOI5Z6V0k6zcUexh0uU3IDqbdudvmWH8zYTo7J2XwR11kp4QgaX1FElmtY
XjSSDKwr+CQZf4tW0ybMozX3o4Rqi73KkgR0IZTEHhnFtz/QMNwcxTAcAMZe81X/
Uhd/A8JGgl4rJELvlQZbLrt6YGqFje5E3xhCg4G5N5qVBciIMZ5tSukLEl+kF+9X
FchFJH0zP2Q5D38fi8h0wAgWBeKeolP3lEdLPgjP7pQuJ1fRxGc5t4xAcNWB1swU
l9Ez72tyi2aKZiK0Gq+LYrKyOPkFRMD+w1M5FNbYy0inhfXoVJ4XudoJ+TGiCte2
nKkUdS3aT7AItZxZqq3TBa8ptv4v3EkKvcGgCjQIJjX0hyvSC0FOc4+1AmJ2MNps
W0+I4+fCjrcquCeHRPbMohjHXmWJyzyJvXXPoLMqdFMOeTkrUV8H2H0HPFgz9kgx
UMXydSOvw0rg9oyA0XTPDwZn3KnNlcJoVhaQqGFHXQZ8X6/c/lgCBQvkES6rFL4R
KghfUdzbDFvky0MtK6T2np5vxoQluFSK/gaRIRVNt2k=
`protect END_PROTECTED
