`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tvTyLdWdKjijReuMDsXmo3a7O9scRiAtI9Z+MuxDAHSxMuKDmJ4hJc/GPqRI2KP7
8cA25Jy6F+dVDGEeUW2VIAcmLRi3+s9DaUl5Z6D0mguMiz1MraYvZ4FtKaCa9bWy
G2cDGs5gjUb//tSU8csIkcmZVXvdUhA8pjXGCbXp5hwrp+al+Ir3fcKmHKi3DMcy
vJc45OIHnUaNSkNtT1XVfpwXKX8rCwoBTFMvjTXumyM14iPW9wZVc9A7SgmXGl4c
4dghMxHPjsLkMrT/EpQWXEIK6lpS1oVeCN722Vy4MyePP/gL+bUl35BrVrtYq0Nf
k71WI8QPhlt5cZCXvodrubSDCk/kCEbSBV+sRgy+A3/aMcbAfPJ7S8Gbgsi7+yG5
kGd4U48g3Ms6p5AAmc6IhdIwJa/erUvh7BtYWfBpj2k0qjZQ06XPZf0524I/FalI
i3WqWsexUlSjXrem928UM1Hx7BCJoVqjrjx31+5fj+/XosvFJxzWAH8Dnkt1sQN/
F2aUt5RdasG4yNYhNjgoqLGb3brcZX925RDnG80i2cClsbhRTmJ0T9nZ4CW1gmex
GC8KEeitBe9QN/lflekUANpeQbcJnYTkgfuYxFUL+sA4wMka3I88Dz8s7OPYr76Z
L0UhdaD6WW5SxrV7T2SWIaV5rS1tLIF2LbtoXDdm7hAVFag+sRJ0+uGP86f2aXoR
6241RaJ5JF7J7w3+qUcOPFBUtdjBaPNZWwwAHI4rCdz7fDTeE4S26ARi4ulGezQs
udL3/l5O/dfD/nwMwfR8xCyK0MkDB7q4518txG5NzdqPvTx9kYccYSyvDQ1Q+4fH
5lEUIpDlIgqjIL+rhttWWwPVAm/GgUsl17q+akfnW+jF5DdCw+UMPQpy0LVGUA4v
nDHhphVfSN4d1hxL1M4tZLseGkPKKHJVtLp6NoLc/9S9E4wnY0L+hC3686LJg2CF
3RGmAbA7+hYTNq7uielMTtfgKd7lZN+C6cQvzaBS8tqqHOz/d9rmEusF1BCYiEcT
X8JkZV+a4IJ8adRWbUGfOnxTrAgkq0oS0AleHWysNLjyDivQhTzAY7D+kc5+RAzX
ljo5yXNwTEk6k5efcfZDdJMGUa7rV1toYOUtKqGPkIrCGKFUxY8lXkKHmG+wp1ZF
A5EABBAUxAuXay0twU3LfBni1YnGsjjRmVljSu9IF3dyyjI+ABFrpilm7tvXVRTY
o7p/+aZirywTA1cX7UEVDmIfu91tdJ3VuBGgx1In6HSgxCYb0FIj74HczNN1PJtO
jEEOn2GKyWLYetm3mH/4pSjWLFvDwXtyQWAE75cLY5vXHICl72V7pGSEmNsnxg5A
x9jd+9k8Td0QsI59OFos0k8ujsbEKrt+pYXR7eEgmNrzJ9cKQCnegKN8qDRx6iIj
QFiqqMQ/Q45CeJM//K6bdzh/6ywAeQMS9EuvJf5BOu1vXXZZ9DYz2VUZyai8juub
5JKj2Lpt/ELT6j7//7CRcXkcVhdBOH8EzlJSLeauAencOMiEDfQj3wlysOStd408
pI92eZ+UiN2mssJc6/LIFjWpuCiX7W6jds1/b3STif5LStpsyKf+YlccOjei1l9+
yIWUoKfIsuclFoHQKrd4QKPJplp/w3bPh8uaHJ4VPNPbnvK8tvM01wSIcNt6NG1/
XFPXdBQUyr8ZUAY8yX9VDFsGsqWk1oMReCsY7vjF9vASVBNOG2XVDyyIam5oZgBw
hhBNfS7IhN12cBDTWipSyiO0LHI/5E9jI+x5PJPNaJEa0cHf7/GRGu/eeUqJ0E5U
XBO3alTmxetGfeEuV18NbiXk1vVqAn5HUAvyk+DthJrUCiyG4vdO/KBSFcrhl/vO
U7PiceQYtVgEsQRvbKBQiaFOvNAOsBEjOrrDvSaJCrqRFd3CRCVWArwLejit/Bse
XyMm3PUp+ftT2JnHvTXYUg0cF5ZwWioWxtzVhy8gO6ou3Fg8AfFYhW06UTV2sxrS
qSw/3ZMbJ1MnT6Wd4dp+0oPATohb3VwebpRzFtMPO6q901Pu0n/knDjRHiG9YJSb
D/rp2o/m4miXHYU6PHvFhnVnnTd7/4j80rn6KWlZOxaH6e0GeyS1gdenYafgYJVm
rZXtBfyeiF9/4SGMKQCz1LJMPCrNdME1o9nbiqbvOOPAhnCeCD6psnMucVo6ph8R
k91gQQ3cDJZWSkPCsovrTRbSWFCluJ/7KQg2bRwAIxehnTKbyu0HW8Dl/hYLyiro
QkSXxoRrKWbH2rX1bnlH2iT90hIxxYKKW2Bu6+GD0ZWLKxwWtcPVxI4OqVSDZJOu
UvO3yu6HmVEhcd3JGcuK27MyowKbLIizcRQRZ+rZAob0xRHBseWCWLkzUJTbwoWq
T+Jt4DwALUKBXk4O1M7WkdNRDoBnMCro9TpJH69QGY5doM2qQ5UkK5lfFdPKvHF/
aVfdWzLgVuVAP/YhXyHnSJxp6I1HmKDxpGLsWYdr8vj1HTQC48goSJ0CrSELIVIL
ILlbrAyS1RCz8MaWilRHd4TvjAcFmDpsoDeSGO+bmnmpuHG1DqKHS4KavCZ+aENe
CgSb677IIp1R9nxTetgzOCvca2rH0GEJzwZWObpJNif5Jd4RopOaYdAvNl4TG8DP
fi8u7mtzglRDdOMBFIgo1ctQlvG+g7rTKkBU/iGl0cPsgvrGb+AhZoLnmwo0QgCs
2pIM8k+AUJIvHh8u9RFD7/QFQBxvFfk5et16ANrqNCIoXOwncvBkC8aNpv9YP86t
J5b+a3aCoBzB1G66Clxme3jwl+iUEQ+OoIE9kGz7rNnfU3LZmH5MzDPR3YtI2Q/g
R8yTO9we1UViGY2nJ3XEwdK+MwqY0lGQq2mtq8ECpLK1a+ZngHM3rDs6N0DyVg+y
WXeW0JYAht1FJt0780e5jTZSh66u9Iu7kATGrT8Fyt1J9t6EJu/D+hOj1huLO3BA
PylySaBd8wwR4kCEoJS58u8MVfCYy+BLVfaPg4yRGIl1pLyWbumQkemZSL57KbRG
hMqq4TpoYNmM1d8ylMcpvwzap+LzD8paVZbmqGQVNVGffkGFGEYVZUI6U+W+IAeK
oMe7UNzqovlwV5t+9WcAcZ3gn9UO+R5v2Ec9q2QqtgxLAeYSC3P9HstV26+Ul0g0
dlllpDwYF33QGJvztWK/0FV3clMtVSuv0AdHuUx/9PbJhboT0fL0QJ9gLs8Y7ppx
WKsjlHIrYn3vPObMLnfZDJ107LZjQ/aM1hPq5xg/3eohO0677cXhzTov3dwe3vWI
ok6nKjVPZi12KFxloWBL0NyTqS0Hv5edFZ5uLN/ybt20PBMT2dDW8gVcPrYMBAe+
XpQzW/X2QTWEMTKrSHPIx99GpivG8cxQC/WBZgqcmqNZdV5ltZRqY0D5wjdZuevp
JBivISYW3cF9lm/8XqSpnsP0PQtHlhNyjORsWjkw7pXqm8/2cDrVQ8xJluQM77jO
n6lDjXwfwcheGz77qRPI1CWZQ1mUWUFfs9ia8SmF8jff+jyySqwjkF7jBN0nyJKe
WIV+geFtxSLUmqQf7pHLKmf7s9wsDJdo2wQ94ODNCWgcI04OQswe6+D27z2l+Mtu
FXTxcqbw0GdV8fx6QkQFkMiWmOJ0dfLa25cFjyxXASUBntl+IkfSfS14ECUYNAGo
3kjqRmwWdrkdA/N6xtGbqXDTk9XTmrFa5ap6d+rXVzvBq7sR/Z5zibtu32eJXCIj
1s1w4b0pjR0nFojln0iATo4n++5tJNl/1EVztAqj34fTwBG+o5ZL3cOAZ/fsmaEo
WFcMLbb0zPkGsmGZXOtEX2vNmjkOdhjMLaHLtupgd7+0F3hh6ayZG3H9Aysk+hUg
qas83Wj5t+nMFcrwFUgL0fozZRLENw/BN/gVa14ZTDTOXNlmibPXFP/vBtiSYJB5
E2JwSOfYRQXij6Mz/RWfsLzP+/fNwZU3xI2DXABb86MFMeLyg/D3vfIBH72LcvS4
FS0uC2OIjqdfbFEutLPi1UpD7/lMC9GQ+pVfuA7tXcupPQvIzpt4m8oOJUpRB9fu
/gL85YrW2pN1dhQM1kECDwiCJtL/BhTAaKPYLKl1FrJbBEc9p57Ur+VXHNq1R72t
Ed/kcQ8dZNw+eTY5JxoYe5yzB7NjZgmlrjBM0XCz3y2pfxe+nTNvRVupAwZCkjh1
NIffpwZASLK10EXq3qBISDHWk0jL15PksCTnpnu9pHFvrFLkXOdeVZOPNLkjasrr
L6z92cVD8kydpr31V3YdgbeY24dZ2pZa1KJBO5GhDWMWHbaGODT49IYIoB5cvC5m
952R6DN2XW0/CfDo7DXP+382dIFxdzDmIN/NoX2L+FFXASKI3grQkR55Ayhn/7jv
JHfZHjv+pfv9bDsOqeysWd8BrQwAOemlz1hqjbcU8q8cmTl1BdAlI1qzSzDnMoPY
Wmrus8bHBDb0Aa3m57UC0do3XN1HF3oLbmMe8NipeazH3SCseCyZpXt4PS4SC8UU
/TphBcq8uO45WplA4IyfBRCg3L4rlyCXlEVdwM7AaBcnwUj7dDDDnbA2WuKm/PD4
hRUpPu9jGhj7sO7SE7acLJMDF8Cfdy7zE+va16UJUKeNja6oEWKMpiQ2ifMj/x9k
129IG1s91Fp4TBoFzHGw9inLvUgOXICzSEd1TkcoeWB/XIOu+ffWvM2L7yyMtTFF
px1RyTjGvKJScOlGVeM2n+Xq//hCOfx/JUQilquUnlN34uZHrkE/mnfl6KgSkidi
bEeCb45yKcW2g7oKO6Yo9i6iTH2mxoycNsqSLwURajjNCKZMPIifeIV3lof8JGcf
mFzaZA6UmQQbqh33kbLyB228wrSQjfwgpW46nZV+9SGBol4iiVKT0KLaEoYJCX3J
Vfn42mow8lJgSiBiIBnvkC4zRQriw3ZEIsr92+N29YqeH4YSTtitAKxyOdKayZDy
Ai1EiG+IeZQ9f580gqJuK4nwFdckJckaJ/6tjYmC6Itvqj4uWxj+xrrpMlFIkIW7
qd5yXe+iofQFfMy8+r6x2xHxuNXqRGiU7+shTb0VVf/SG/5nCNqCKvD8jC03l8vo
3uxxvavcKn/hJ00a/wYnfsrWtb0UMAqgWvzGMwMfgB9Pesrt7CmejGYmeWhXVLAS
Q/OUyZSfIUdvr3YtRM95BxUiTfuI9g536MH41SHtkVMvrM1435cgaYjZehOUmNOa
8HmCqT4uGFEjI+jQSInH5VxvWaBz4tJIzR2JW6gsLaCdI2f/78Tw94LLBGNo93WQ
2YjoWqyyL8UqYO3hziBVp+6Peaq3q3rvnwBIQIL7hrhQTVHkgAvYDUw+78H4ENn2
jea62rOSqUf8OHQx2ZG79L2XvLUs/7R9DUeXeIPmhJ5aSpT13Y79o/QgGDI1JtI+
RcrO1LnK2Dlb256DAgK45VRXKDlOAV+rdWp519H+iPiteV3qO11qkzSUZE9QQY6C
y+mQEePKrsjdFFgXE3hFYPE6VFtok9qveaOLfYFQCfZSJf9m38Y83/2iO0MwSIAx
M0ZTzjMsFt/p9ZYovEe6MZPjuzfeL65i7PrSX2W7cdr2+pkVg9Qvy1yiOJemBeJC
n4+Pv9ROvTXQbuHBmT3rlVUxPExzZuQrcYxlq71n2hiOciVrG+K+hymCcwm46mzN
K51e6xQUFtLjF9bm+tanMvu1nQZafjLiodddTVRB4xfOz70qBwh1rRZkAWBstWHG
zeZqyR+aerNATOx+IhGUBRS7PAUBmxag+APpggCXRZy5qMqiUxeqoAp7RpCHnxl0
bBw34+mgNXPw+goF4EuzLusXBmhLWwKcZLjhl2IGpM6HRBFvGw3QAx42DSi8k/2f
HDowUzyyeZ03FwSybRsAksU67oBAo/VYKjmFeA9m9rij/XzqsnJeloyBLUnAr5Yw
xmfGuNi0LH79KA5LRK7VJeZZ50iW9btUR3QgXnvaDOOglL0+hFVsO88HQhisBA7Y
Bge4nankY0t1IBasrIUobkejzF8SuNl9/kIKfLXZW8H4rb9YTKpsvnd7CTVyll1v
auJbeRQaUTke2taHvbAzD6e6CX2bEi/PB4H4G2BoCXE=
`protect END_PROTECTED
