`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+AVSkvMN9xNbrDby/39slcVhjDhhB6tNGGay9u9rZPp3o+BjgKbhOKJ5zrL33Jku
2Y5AHmoM0M7KTsCwsQT/0JZwk5eUTGA7wIdTPKO31n0K4+u/ld0HrS4XPXCtyqhx
4XFh5e9/DaqpMXzI96me0aG5IC4PKpv3/8B2EYa7KgyL9QpyLIJORn3B0/JzZztB
NqZS9Y5EPTX7pGuw7isfAeDBzeotDF12XDLu9v+8ukuI7EV3ts35Pbu/c9bhk994
o2i1vDcmOMFN01/gHoxYboB9VpwBQOP9JYPGgrqXRkvUJ3UEdcv680kGvnj7MOEl
RY7uXJ2P4Dfqa8KYAeA2Gyq6/Xeq0zR/WqIO4ws/Fw/uwUUgjnlM+1QwxRmhff7F
iIZbgDIUJX5mABS/eppxPkpqr+V1X9xwxSS0Z5rQRYf36jVJ8vZAIbHytPQCjf2E
4mbguC2Wio8P4noTurx6jTx46Qt1CpzreRHZLiWStp8LPQFGmOzdj02PGYGAbqZ3
X/5jUsqjRNoNFdotmvJeca0peNJzbqfRnkD/T5zHWzU2H8Q6+HN0CIwvbraIUil+
4vCLBsNLIlvF77Zz3L45JtY+JQUBSMmFmHxcYLRLXzJnCFAyrT2wx2J3vIOPC7gN
/+6uef7qFCLE1EcJqPSBGcJDRh3ahYBlkoLxznJd8oQ2aSmLIdtLoDUzN4coTCjx
z0ihSZRk7xRMm27YF9e4R0T+WWIAepv+6UDne+XQ9KOzv0fnpLPb0jlBUDWluUOz
KOLrq3uIl5Pf5NMmXTGPzmmz5qXPxXSWoO4XwNlJ/S1ntUbt3zUHli7d+jPzW1lc
0pIOHMb4A3SEqNQpOqkhmSNt8orQWwbrRUyvEIrhmEXXtRBKOyTRnEnjJv1C38ay
UPm/UCApzVdp6dPonQihBDOlH8eXc6OL9SeHamOeoiTxA5h9q2XSk5HjfZ+sbc8m
iPtPv4OsxzSObVE/VbC1CfBIBrGXb+cFFI5T6Hf8anF/RoOmvHQIYjWJOwFze2OA
6otrJDHB2L2lJSejM+/aOFWRjQAVhdJyOvsMxdiPMjye2AypMuw3+s2TCiLEAblj
gqcEptFJ+BoRaKWA2qsCtqh9A2kcC3v9R+Xjno634aaJ8e+f2HrOF26Z/2MH2s8T
4afadCUOnZGE0j4OuTxmY13yEmM2hlAI4b1SyQdTM1cJ91jta4sI9te1JExK3MOJ
nnzNNdetZMyAGK1ls0514WP/6QMLLv05TMgd9Ha/SxLM7dvsF0jxK2xAL55aK3eu
EowJBQuoF+IKJfKiMYHBtnOyEUN4uznxEtrFd/68V73zrvFsAkWL0bFUOB8FM+5t
Ay2Jl+M9hTwIm+wLLNe0AscL+d1rrBUs7ZZC2cwGgew0QOAy5Z4EWMNYiAa/gM4J
u/IHzJIm8pX9Z6fCr0kRrwrCwXb8ph8jm7w9XKkoEV2XldeuxstbeN+xnWBug5Rh
jlLwPq+SWHCEUWvsO0ohskqZ3sv12e7wPFt8uiJ5LZbt0GIajGz4CZ7KtBmgXTEi
WltOflvHI2QU4i82/P2msksuwff/uHkLMKHxZht0yK4cIGG+l5jB7ZNw+CUUa3q/
TASHbDa+tmGIKwtglHg2OzVFQ/PanExZA6RXH1oFAK4RiLWQdFO18BoLLhVzJKNK
evn7FE4m29P985T3Hhy0lePKwo+din/2jen0FnrqVm0YnvpNIXRwBSLBL3dh0k/+
oqea8QjH0EMZS8D2Ppdrz6x63Q9E2NJo0JJbQ0M1ZGGk+S18MN9VsJF8TlZsairL
R77S8yoyKUb7SBPDJ5IYVTKle1TKQCu+4QT3QGcKvncikh6jYa5BPm0nqK54h9uv
qLzmvhcQ2NS06sW+PJ8uf85/xrxZ270FYBaFHVJNpIQEMlJW1qmk4GiV5It3YJKs
pGEPOw+mcgpS0BB8I7DkhdmE6DSyFG/6oGZP0vFOPebUnDWGV7SbvB0OmPoc0KFU
6LN/lBvHt7W3EZs0g6eYNGBEX0Lz7uxfK2uhhxSg3qhEYqMv8nV8IKG5v419pSja
l7cv45eqG4o2DLruuGQhiEvfbLesUSHvKoJodtmWSnyW1c+ReLGpbYxT3Aajl5ET
LGm5t5/Y1+2ZKPEeAIGm0Vv5WxJfEWes0dedZX81pOfJ+/gx3sBRV3YLc+yhM0kH
6u8BWOp/EAKEONfUpVkAv7A9DsHy+xy0vIfMNnhgAidhxvm4SXadyR2xONaMqi6V
jfeDlQbIXyiT+slrkkUX4Q==
`protect END_PROTECTED
